
module FIFO_DEPTH_P25_WIDTH16 ( clk, reset, data_in, put, get, data_out, empty, 
        full, fillcount );
  input [15:0] data_in;
  output [15:0] data_out;
  output [5:0] fillcount;
  input clk, reset, put, get;
  output empty, full;
  wire   n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n50, n51, n52, n53, n55, n56, n57,
         n58, n66, n67, n68, n69, n70, n77, n78, n79, n80, n81, n82, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n54, n59, n60, n61, n62, n63,
         n64, n65, n71, n72, n73, n74, n75, n76, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n119,
         n137, n155, n173, n191, n209, n227, n245, n263, n280, n297, n314,
         n331, n348, n365, n382, n400, n417, n434, n451, n468, n485, n502,
         n519, n537, n554, n571, n588, n605, n622, n639, n666, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350;
  wire   [4:0] wr_ptr;
  wire   [511:0] fifo_array;
  wire   [5:2] add_45_carry;
  wire   [4:2] r308_carry;
  wire   [4:2] r307_carry;

  DFFPOSX1 full_reg ( .D(n1239), .CLK(clk), .Q(full) );
  DFFPOSX1 fillcount_reg_5_ ( .D(n1238), .CLK(clk), .Q(fillcount[5]) );
  DFFPOSX1 empty_reg ( .D(n1237), .CLK(clk), .Q(empty) );
  DFFPOSX1 wr_ptr_reg_0_ ( .D(n1231), .CLK(clk), .Q(wr_ptr[0]) );
  DFFPOSX1 wr_ptr_reg_1_ ( .D(n1230), .CLK(clk), .Q(wr_ptr[1]) );
  DFFPOSX1 wr_ptr_reg_2_ ( .D(n1229), .CLK(clk), .Q(wr_ptr[2]) );
  DFFPOSX1 wr_ptr_reg_3_ ( .D(n1228), .CLK(clk), .Q(wr_ptr[3]) );
  DFFPOSX1 wr_ptr_reg_4_ ( .D(n1227), .CLK(clk), .Q(wr_ptr[4]) );
  DFFPOSX1 data_out_reg_0_ ( .D(n2320), .CLK(clk), .Q(data_out[0]) );
  DFFPOSX1 data_out_reg_1_ ( .D(n2321), .CLK(clk), .Q(data_out[1]) );
  DFFPOSX1 data_out_reg_2_ ( .D(n2322), .CLK(clk), .Q(data_out[2]) );
  DFFPOSX1 data_out_reg_3_ ( .D(n2323), .CLK(clk), .Q(data_out[3]) );
  DFFPOSX1 data_out_reg_4_ ( .D(n2324), .CLK(clk), .Q(data_out[4]) );
  DFFPOSX1 data_out_reg_5_ ( .D(n2325), .CLK(clk), .Q(data_out[5]) );
  DFFPOSX1 data_out_reg_6_ ( .D(n2326), .CLK(clk), .Q(data_out[6]) );
  DFFPOSX1 data_out_reg_7_ ( .D(n2327), .CLK(clk), .Q(data_out[7]) );
  DFFPOSX1 data_out_reg_8_ ( .D(n2328), .CLK(clk), .Q(data_out[8]) );
  DFFPOSX1 data_out_reg_9_ ( .D(n2329), .CLK(clk), .Q(data_out[9]) );
  DFFPOSX1 data_out_reg_10_ ( .D(n2330), .CLK(clk), .Q(data_out[10]) );
  DFFPOSX1 data_out_reg_11_ ( .D(n2331), .CLK(clk), .Q(data_out[11]) );
  DFFPOSX1 data_out_reg_12_ ( .D(n2332), .CLK(clk), .Q(data_out[12]) );
  DFFPOSX1 data_out_reg_13_ ( .D(n2333), .CLK(clk), .Q(data_out[13]) );
  DFFPOSX1 data_out_reg_14_ ( .D(n2334), .CLK(clk), .Q(data_out[14]) );
  DFFPOSX1 data_out_reg_15_ ( .D(n2335), .CLK(clk), .Q(data_out[15]) );
  DFFPOSX1 rd_ptr_reg_0_ ( .D(n2336), .CLK(clk), .Q(n19) );
  DFFPOSX1 rd_ptr_reg_1_ ( .D(n2337), .CLK(clk), .Q(n20) );
  DFFPOSX1 rd_ptr_reg_2_ ( .D(n2338), .CLK(clk), .Q(n21) );
  DFFPOSX1 rd_ptr_reg_3_ ( .D(n2339), .CLK(clk), .Q(n22) );
  DFFPOSX1 rd_ptr_reg_4_ ( .D(n2340), .CLK(clk), .Q(n23) );
  DFFPOSX1 fillcount_reg_0_ ( .D(n1236), .CLK(clk), .Q(fillcount[0]) );
  DFFPOSX1 fillcount_reg_4_ ( .D(n1232), .CLK(clk), .Q(fillcount[4]) );
  DFFPOSX1 fillcount_reg_1_ ( .D(n1235), .CLK(clk), .Q(fillcount[1]) );
  DFFPOSX1 fillcount_reg_2_ ( .D(n1234), .CLK(clk), .Q(fillcount[2]) );
  DFFPOSX1 fillcount_reg_3_ ( .D(n1233), .CLK(clk), .Q(fillcount[3]) );
  DFFPOSX1 fifo_array_reg_31__15_ ( .D(n1226), .CLK(clk), .Q(fifo_array[511])
         );
  DFFPOSX1 fifo_array_reg_31__14_ ( .D(n1225), .CLK(clk), .Q(fifo_array[510])
         );
  DFFPOSX1 fifo_array_reg_31__13_ ( .D(n1224), .CLK(clk), .Q(fifo_array[509])
         );
  DFFPOSX1 fifo_array_reg_31__12_ ( .D(n1223), .CLK(clk), .Q(fifo_array[508])
         );
  DFFPOSX1 fifo_array_reg_31__11_ ( .D(n1222), .CLK(clk), .Q(fifo_array[507])
         );
  DFFPOSX1 fifo_array_reg_31__10_ ( .D(n1221), .CLK(clk), .Q(fifo_array[506])
         );
  DFFPOSX1 fifo_array_reg_31__9_ ( .D(n1220), .CLK(clk), .Q(fifo_array[505])
         );
  DFFPOSX1 fifo_array_reg_31__8_ ( .D(n1219), .CLK(clk), .Q(fifo_array[504])
         );
  DFFPOSX1 fifo_array_reg_31__7_ ( .D(n1218), .CLK(clk), .Q(fifo_array[503])
         );
  DFFPOSX1 fifo_array_reg_31__6_ ( .D(n1217), .CLK(clk), .Q(fifo_array[502])
         );
  DFFPOSX1 fifo_array_reg_31__5_ ( .D(n1216), .CLK(clk), .Q(fifo_array[501])
         );
  DFFPOSX1 fifo_array_reg_31__4_ ( .D(n1215), .CLK(clk), .Q(fifo_array[500])
         );
  DFFPOSX1 fifo_array_reg_31__3_ ( .D(n1214), .CLK(clk), .Q(fifo_array[499])
         );
  DFFPOSX1 fifo_array_reg_31__2_ ( .D(n1213), .CLK(clk), .Q(fifo_array[498])
         );
  DFFPOSX1 fifo_array_reg_31__1_ ( .D(n1212), .CLK(clk), .Q(fifo_array[497])
         );
  DFFPOSX1 fifo_array_reg_31__0_ ( .D(n1211), .CLK(clk), .Q(fifo_array[496])
         );
  DFFPOSX1 fifo_array_reg_30__15_ ( .D(n1210), .CLK(clk), .Q(fifo_array[495])
         );
  DFFPOSX1 fifo_array_reg_30__14_ ( .D(n1209), .CLK(clk), .Q(fifo_array[494])
         );
  DFFPOSX1 fifo_array_reg_30__13_ ( .D(n1208), .CLK(clk), .Q(fifo_array[493])
         );
  DFFPOSX1 fifo_array_reg_30__12_ ( .D(n1207), .CLK(clk), .Q(fifo_array[492])
         );
  DFFPOSX1 fifo_array_reg_30__11_ ( .D(n1206), .CLK(clk), .Q(fifo_array[491])
         );
  DFFPOSX1 fifo_array_reg_30__10_ ( .D(n1205), .CLK(clk), .Q(fifo_array[490])
         );
  DFFPOSX1 fifo_array_reg_30__9_ ( .D(n1204), .CLK(clk), .Q(fifo_array[489])
         );
  DFFPOSX1 fifo_array_reg_30__8_ ( .D(n1203), .CLK(clk), .Q(fifo_array[488])
         );
  DFFPOSX1 fifo_array_reg_30__7_ ( .D(n1202), .CLK(clk), .Q(fifo_array[487])
         );
  DFFPOSX1 fifo_array_reg_30__6_ ( .D(n1201), .CLK(clk), .Q(fifo_array[486])
         );
  DFFPOSX1 fifo_array_reg_30__5_ ( .D(n1200), .CLK(clk), .Q(fifo_array[485])
         );
  DFFPOSX1 fifo_array_reg_30__4_ ( .D(n1199), .CLK(clk), .Q(fifo_array[484])
         );
  DFFPOSX1 fifo_array_reg_30__3_ ( .D(n1198), .CLK(clk), .Q(fifo_array[483])
         );
  DFFPOSX1 fifo_array_reg_30__2_ ( .D(n1197), .CLK(clk), .Q(fifo_array[482])
         );
  DFFPOSX1 fifo_array_reg_30__1_ ( .D(n1196), .CLK(clk), .Q(fifo_array[481])
         );
  DFFPOSX1 fifo_array_reg_30__0_ ( .D(n1195), .CLK(clk), .Q(fifo_array[480])
         );
  DFFPOSX1 fifo_array_reg_29__15_ ( .D(n1194), .CLK(clk), .Q(fifo_array[479])
         );
  DFFPOSX1 fifo_array_reg_29__14_ ( .D(n1193), .CLK(clk), .Q(fifo_array[478])
         );
  DFFPOSX1 fifo_array_reg_29__13_ ( .D(n1192), .CLK(clk), .Q(fifo_array[477])
         );
  DFFPOSX1 fifo_array_reg_29__12_ ( .D(n1191), .CLK(clk), .Q(fifo_array[476])
         );
  DFFPOSX1 fifo_array_reg_29__11_ ( .D(n1190), .CLK(clk), .Q(fifo_array[475])
         );
  DFFPOSX1 fifo_array_reg_29__10_ ( .D(n1189), .CLK(clk), .Q(fifo_array[474])
         );
  DFFPOSX1 fifo_array_reg_29__9_ ( .D(n1188), .CLK(clk), .Q(fifo_array[473])
         );
  DFFPOSX1 fifo_array_reg_29__8_ ( .D(n1187), .CLK(clk), .Q(fifo_array[472])
         );
  DFFPOSX1 fifo_array_reg_29__7_ ( .D(n1186), .CLK(clk), .Q(fifo_array[471])
         );
  DFFPOSX1 fifo_array_reg_29__6_ ( .D(n1185), .CLK(clk), .Q(fifo_array[470])
         );
  DFFPOSX1 fifo_array_reg_29__5_ ( .D(n1184), .CLK(clk), .Q(fifo_array[469])
         );
  DFFPOSX1 fifo_array_reg_29__4_ ( .D(n1183), .CLK(clk), .Q(fifo_array[468])
         );
  DFFPOSX1 fifo_array_reg_29__3_ ( .D(n1182), .CLK(clk), .Q(fifo_array[467])
         );
  DFFPOSX1 fifo_array_reg_29__2_ ( .D(n1181), .CLK(clk), .Q(fifo_array[466])
         );
  DFFPOSX1 fifo_array_reg_29__1_ ( .D(n1180), .CLK(clk), .Q(fifo_array[465])
         );
  DFFPOSX1 fifo_array_reg_29__0_ ( .D(n1179), .CLK(clk), .Q(fifo_array[464])
         );
  DFFPOSX1 fifo_array_reg_28__15_ ( .D(n1178), .CLK(clk), .Q(fifo_array[463])
         );
  DFFPOSX1 fifo_array_reg_28__14_ ( .D(n1177), .CLK(clk), .Q(fifo_array[462])
         );
  DFFPOSX1 fifo_array_reg_28__13_ ( .D(n1176), .CLK(clk), .Q(fifo_array[461])
         );
  DFFPOSX1 fifo_array_reg_28__12_ ( .D(n1175), .CLK(clk), .Q(fifo_array[460])
         );
  DFFPOSX1 fifo_array_reg_28__11_ ( .D(n1174), .CLK(clk), .Q(fifo_array[459])
         );
  DFFPOSX1 fifo_array_reg_28__10_ ( .D(n1173), .CLK(clk), .Q(fifo_array[458])
         );
  DFFPOSX1 fifo_array_reg_28__9_ ( .D(n1172), .CLK(clk), .Q(fifo_array[457])
         );
  DFFPOSX1 fifo_array_reg_28__8_ ( .D(n1171), .CLK(clk), .Q(fifo_array[456])
         );
  DFFPOSX1 fifo_array_reg_28__7_ ( .D(n1170), .CLK(clk), .Q(fifo_array[455])
         );
  DFFPOSX1 fifo_array_reg_28__6_ ( .D(n1169), .CLK(clk), .Q(fifo_array[454])
         );
  DFFPOSX1 fifo_array_reg_28__5_ ( .D(n1168), .CLK(clk), .Q(fifo_array[453])
         );
  DFFPOSX1 fifo_array_reg_28__4_ ( .D(n1167), .CLK(clk), .Q(fifo_array[452])
         );
  DFFPOSX1 fifo_array_reg_28__3_ ( .D(n1166), .CLK(clk), .Q(fifo_array[451])
         );
  DFFPOSX1 fifo_array_reg_28__2_ ( .D(n1165), .CLK(clk), .Q(fifo_array[450])
         );
  DFFPOSX1 fifo_array_reg_28__1_ ( .D(n1164), .CLK(clk), .Q(fifo_array[449])
         );
  DFFPOSX1 fifo_array_reg_28__0_ ( .D(n1163), .CLK(clk), .Q(fifo_array[448])
         );
  DFFPOSX1 fifo_array_reg_27__15_ ( .D(n1162), .CLK(clk), .Q(fifo_array[447])
         );
  DFFPOSX1 fifo_array_reg_27__14_ ( .D(n1161), .CLK(clk), .Q(fifo_array[446])
         );
  DFFPOSX1 fifo_array_reg_27__13_ ( .D(n1160), .CLK(clk), .Q(fifo_array[445])
         );
  DFFPOSX1 fifo_array_reg_27__12_ ( .D(n1159), .CLK(clk), .Q(fifo_array[444])
         );
  DFFPOSX1 fifo_array_reg_27__11_ ( .D(n1158), .CLK(clk), .Q(fifo_array[443])
         );
  DFFPOSX1 fifo_array_reg_27__10_ ( .D(n1157), .CLK(clk), .Q(fifo_array[442])
         );
  DFFPOSX1 fifo_array_reg_27__9_ ( .D(n1156), .CLK(clk), .Q(fifo_array[441])
         );
  DFFPOSX1 fifo_array_reg_27__8_ ( .D(n1155), .CLK(clk), .Q(fifo_array[440])
         );
  DFFPOSX1 fifo_array_reg_27__7_ ( .D(n1154), .CLK(clk), .Q(fifo_array[439])
         );
  DFFPOSX1 fifo_array_reg_27__6_ ( .D(n1153), .CLK(clk), .Q(fifo_array[438])
         );
  DFFPOSX1 fifo_array_reg_27__5_ ( .D(n1152), .CLK(clk), .Q(fifo_array[437])
         );
  DFFPOSX1 fifo_array_reg_27__4_ ( .D(n1151), .CLK(clk), .Q(fifo_array[436])
         );
  DFFPOSX1 fifo_array_reg_27__3_ ( .D(n1150), .CLK(clk), .Q(fifo_array[435])
         );
  DFFPOSX1 fifo_array_reg_27__2_ ( .D(n1149), .CLK(clk), .Q(fifo_array[434])
         );
  DFFPOSX1 fifo_array_reg_27__1_ ( .D(n1148), .CLK(clk), .Q(fifo_array[433])
         );
  DFFPOSX1 fifo_array_reg_27__0_ ( .D(n1147), .CLK(clk), .Q(fifo_array[432])
         );
  DFFPOSX1 fifo_array_reg_26__15_ ( .D(n1146), .CLK(clk), .Q(fifo_array[431])
         );
  DFFPOSX1 fifo_array_reg_26__14_ ( .D(n1145), .CLK(clk), .Q(fifo_array[430])
         );
  DFFPOSX1 fifo_array_reg_26__13_ ( .D(n1144), .CLK(clk), .Q(fifo_array[429])
         );
  DFFPOSX1 fifo_array_reg_26__12_ ( .D(n1143), .CLK(clk), .Q(fifo_array[428])
         );
  DFFPOSX1 fifo_array_reg_26__11_ ( .D(n1142), .CLK(clk), .Q(fifo_array[427])
         );
  DFFPOSX1 fifo_array_reg_26__10_ ( .D(n1141), .CLK(clk), .Q(fifo_array[426])
         );
  DFFPOSX1 fifo_array_reg_26__9_ ( .D(n1140), .CLK(clk), .Q(fifo_array[425])
         );
  DFFPOSX1 fifo_array_reg_26__8_ ( .D(n1139), .CLK(clk), .Q(fifo_array[424])
         );
  DFFPOSX1 fifo_array_reg_26__7_ ( .D(n1138), .CLK(clk), .Q(fifo_array[423])
         );
  DFFPOSX1 fifo_array_reg_26__6_ ( .D(n1137), .CLK(clk), .Q(fifo_array[422])
         );
  DFFPOSX1 fifo_array_reg_26__5_ ( .D(n1136), .CLK(clk), .Q(fifo_array[421])
         );
  DFFPOSX1 fifo_array_reg_26__4_ ( .D(n1135), .CLK(clk), .Q(fifo_array[420])
         );
  DFFPOSX1 fifo_array_reg_26__3_ ( .D(n1134), .CLK(clk), .Q(fifo_array[419])
         );
  DFFPOSX1 fifo_array_reg_26__2_ ( .D(n1133), .CLK(clk), .Q(fifo_array[418])
         );
  DFFPOSX1 fifo_array_reg_26__1_ ( .D(n1132), .CLK(clk), .Q(fifo_array[417])
         );
  DFFPOSX1 fifo_array_reg_26__0_ ( .D(n1131), .CLK(clk), .Q(fifo_array[416])
         );
  DFFPOSX1 fifo_array_reg_25__15_ ( .D(n1130), .CLK(clk), .Q(fifo_array[415])
         );
  DFFPOSX1 fifo_array_reg_25__14_ ( .D(n1129), .CLK(clk), .Q(fifo_array[414])
         );
  DFFPOSX1 fifo_array_reg_25__13_ ( .D(n1128), .CLK(clk), .Q(fifo_array[413])
         );
  DFFPOSX1 fifo_array_reg_25__12_ ( .D(n1127), .CLK(clk), .Q(fifo_array[412])
         );
  DFFPOSX1 fifo_array_reg_25__11_ ( .D(n1126), .CLK(clk), .Q(fifo_array[411])
         );
  DFFPOSX1 fifo_array_reg_25__10_ ( .D(n1125), .CLK(clk), .Q(fifo_array[410])
         );
  DFFPOSX1 fifo_array_reg_25__9_ ( .D(n1124), .CLK(clk), .Q(fifo_array[409])
         );
  DFFPOSX1 fifo_array_reg_25__8_ ( .D(n1123), .CLK(clk), .Q(fifo_array[408])
         );
  DFFPOSX1 fifo_array_reg_25__7_ ( .D(n1122), .CLK(clk), .Q(fifo_array[407])
         );
  DFFPOSX1 fifo_array_reg_25__6_ ( .D(n1121), .CLK(clk), .Q(fifo_array[406])
         );
  DFFPOSX1 fifo_array_reg_25__5_ ( .D(n1120), .CLK(clk), .Q(fifo_array[405])
         );
  DFFPOSX1 fifo_array_reg_25__4_ ( .D(n1119), .CLK(clk), .Q(fifo_array[404])
         );
  DFFPOSX1 fifo_array_reg_25__3_ ( .D(n1118), .CLK(clk), .Q(fifo_array[403])
         );
  DFFPOSX1 fifo_array_reg_25__2_ ( .D(n1117), .CLK(clk), .Q(fifo_array[402])
         );
  DFFPOSX1 fifo_array_reg_25__1_ ( .D(n1116), .CLK(clk), .Q(fifo_array[401])
         );
  DFFPOSX1 fifo_array_reg_25__0_ ( .D(n1115), .CLK(clk), .Q(fifo_array[400])
         );
  DFFPOSX1 fifo_array_reg_24__15_ ( .D(n1114), .CLK(clk), .Q(fifo_array[399])
         );
  DFFPOSX1 fifo_array_reg_24__14_ ( .D(n1113), .CLK(clk), .Q(fifo_array[398])
         );
  DFFPOSX1 fifo_array_reg_24__13_ ( .D(n1112), .CLK(clk), .Q(fifo_array[397])
         );
  DFFPOSX1 fifo_array_reg_24__12_ ( .D(n1111), .CLK(clk), .Q(fifo_array[396])
         );
  DFFPOSX1 fifo_array_reg_24__11_ ( .D(n1110), .CLK(clk), .Q(fifo_array[395])
         );
  DFFPOSX1 fifo_array_reg_24__10_ ( .D(n1109), .CLK(clk), .Q(fifo_array[394])
         );
  DFFPOSX1 fifo_array_reg_24__9_ ( .D(n1108), .CLK(clk), .Q(fifo_array[393])
         );
  DFFPOSX1 fifo_array_reg_24__8_ ( .D(n1107), .CLK(clk), .Q(fifo_array[392])
         );
  DFFPOSX1 fifo_array_reg_24__7_ ( .D(n1106), .CLK(clk), .Q(fifo_array[391])
         );
  DFFPOSX1 fifo_array_reg_24__6_ ( .D(n1105), .CLK(clk), .Q(fifo_array[390])
         );
  DFFPOSX1 fifo_array_reg_24__5_ ( .D(n1104), .CLK(clk), .Q(fifo_array[389])
         );
  DFFPOSX1 fifo_array_reg_24__4_ ( .D(n1103), .CLK(clk), .Q(fifo_array[388])
         );
  DFFPOSX1 fifo_array_reg_24__3_ ( .D(n1102), .CLK(clk), .Q(fifo_array[387])
         );
  DFFPOSX1 fifo_array_reg_24__2_ ( .D(n1101), .CLK(clk), .Q(fifo_array[386])
         );
  DFFPOSX1 fifo_array_reg_24__1_ ( .D(n1100), .CLK(clk), .Q(fifo_array[385])
         );
  DFFPOSX1 fifo_array_reg_24__0_ ( .D(n1099), .CLK(clk), .Q(fifo_array[384])
         );
  DFFPOSX1 fifo_array_reg_23__15_ ( .D(n1098), .CLK(clk), .Q(fifo_array[383])
         );
  DFFPOSX1 fifo_array_reg_23__14_ ( .D(n1097), .CLK(clk), .Q(fifo_array[382])
         );
  DFFPOSX1 fifo_array_reg_23__13_ ( .D(n1096), .CLK(clk), .Q(fifo_array[381])
         );
  DFFPOSX1 fifo_array_reg_23__12_ ( .D(n1095), .CLK(clk), .Q(fifo_array[380])
         );
  DFFPOSX1 fifo_array_reg_23__11_ ( .D(n1094), .CLK(clk), .Q(fifo_array[379])
         );
  DFFPOSX1 fifo_array_reg_23__10_ ( .D(n1093), .CLK(clk), .Q(fifo_array[378])
         );
  DFFPOSX1 fifo_array_reg_23__9_ ( .D(n1092), .CLK(clk), .Q(fifo_array[377])
         );
  DFFPOSX1 fifo_array_reg_23__8_ ( .D(n1091), .CLK(clk), .Q(fifo_array[376])
         );
  DFFPOSX1 fifo_array_reg_23__7_ ( .D(n1090), .CLK(clk), .Q(fifo_array[375])
         );
  DFFPOSX1 fifo_array_reg_23__6_ ( .D(n1089), .CLK(clk), .Q(fifo_array[374])
         );
  DFFPOSX1 fifo_array_reg_23__5_ ( .D(n1088), .CLK(clk), .Q(fifo_array[373])
         );
  DFFPOSX1 fifo_array_reg_23__4_ ( .D(n1087), .CLK(clk), .Q(fifo_array[372])
         );
  DFFPOSX1 fifo_array_reg_23__3_ ( .D(n1086), .CLK(clk), .Q(fifo_array[371])
         );
  DFFPOSX1 fifo_array_reg_23__2_ ( .D(n1085), .CLK(clk), .Q(fifo_array[370])
         );
  DFFPOSX1 fifo_array_reg_23__1_ ( .D(n1084), .CLK(clk), .Q(fifo_array[369])
         );
  DFFPOSX1 fifo_array_reg_23__0_ ( .D(n1083), .CLK(clk), .Q(fifo_array[368])
         );
  DFFPOSX1 fifo_array_reg_22__15_ ( .D(n1082), .CLK(clk), .Q(fifo_array[367])
         );
  DFFPOSX1 fifo_array_reg_22__14_ ( .D(n1081), .CLK(clk), .Q(fifo_array[366])
         );
  DFFPOSX1 fifo_array_reg_22__13_ ( .D(n1080), .CLK(clk), .Q(fifo_array[365])
         );
  DFFPOSX1 fifo_array_reg_22__12_ ( .D(n1079), .CLK(clk), .Q(fifo_array[364])
         );
  DFFPOSX1 fifo_array_reg_22__11_ ( .D(n1078), .CLK(clk), .Q(fifo_array[363])
         );
  DFFPOSX1 fifo_array_reg_22__10_ ( .D(n1077), .CLK(clk), .Q(fifo_array[362])
         );
  DFFPOSX1 fifo_array_reg_22__9_ ( .D(n1076), .CLK(clk), .Q(fifo_array[361])
         );
  DFFPOSX1 fifo_array_reg_22__8_ ( .D(n1075), .CLK(clk), .Q(fifo_array[360])
         );
  DFFPOSX1 fifo_array_reg_22__7_ ( .D(n1074), .CLK(clk), .Q(fifo_array[359])
         );
  DFFPOSX1 fifo_array_reg_22__6_ ( .D(n1073), .CLK(clk), .Q(fifo_array[358])
         );
  DFFPOSX1 fifo_array_reg_22__5_ ( .D(n1072), .CLK(clk), .Q(fifo_array[357])
         );
  DFFPOSX1 fifo_array_reg_22__4_ ( .D(n1071), .CLK(clk), .Q(fifo_array[356])
         );
  DFFPOSX1 fifo_array_reg_22__3_ ( .D(n1070), .CLK(clk), .Q(fifo_array[355])
         );
  DFFPOSX1 fifo_array_reg_22__2_ ( .D(n1069), .CLK(clk), .Q(fifo_array[354])
         );
  DFFPOSX1 fifo_array_reg_22__1_ ( .D(n1068), .CLK(clk), .Q(fifo_array[353])
         );
  DFFPOSX1 fifo_array_reg_22__0_ ( .D(n1067), .CLK(clk), .Q(fifo_array[352])
         );
  DFFPOSX1 fifo_array_reg_21__15_ ( .D(n1066), .CLK(clk), .Q(fifo_array[351])
         );
  DFFPOSX1 fifo_array_reg_21__14_ ( .D(n1065), .CLK(clk), .Q(fifo_array[350])
         );
  DFFPOSX1 fifo_array_reg_21__13_ ( .D(n1064), .CLK(clk), .Q(fifo_array[349])
         );
  DFFPOSX1 fifo_array_reg_21__12_ ( .D(n1063), .CLK(clk), .Q(fifo_array[348])
         );
  DFFPOSX1 fifo_array_reg_21__11_ ( .D(n1062), .CLK(clk), .Q(fifo_array[347])
         );
  DFFPOSX1 fifo_array_reg_21__10_ ( .D(n1061), .CLK(clk), .Q(fifo_array[346])
         );
  DFFPOSX1 fifo_array_reg_21__9_ ( .D(n1060), .CLK(clk), .Q(fifo_array[345])
         );
  DFFPOSX1 fifo_array_reg_21__8_ ( .D(n1059), .CLK(clk), .Q(fifo_array[344])
         );
  DFFPOSX1 fifo_array_reg_21__7_ ( .D(n1058), .CLK(clk), .Q(fifo_array[343])
         );
  DFFPOSX1 fifo_array_reg_21__6_ ( .D(n1057), .CLK(clk), .Q(fifo_array[342])
         );
  DFFPOSX1 fifo_array_reg_21__5_ ( .D(n1056), .CLK(clk), .Q(fifo_array[341])
         );
  DFFPOSX1 fifo_array_reg_21__4_ ( .D(n1055), .CLK(clk), .Q(fifo_array[340])
         );
  DFFPOSX1 fifo_array_reg_21__3_ ( .D(n1054), .CLK(clk), .Q(fifo_array[339])
         );
  DFFPOSX1 fifo_array_reg_21__2_ ( .D(n1053), .CLK(clk), .Q(fifo_array[338])
         );
  DFFPOSX1 fifo_array_reg_21__1_ ( .D(n1052), .CLK(clk), .Q(fifo_array[337])
         );
  DFFPOSX1 fifo_array_reg_21__0_ ( .D(n1051), .CLK(clk), .Q(fifo_array[336])
         );
  DFFPOSX1 fifo_array_reg_20__15_ ( .D(n1050), .CLK(clk), .Q(fifo_array[335])
         );
  DFFPOSX1 fifo_array_reg_20__14_ ( .D(n1049), .CLK(clk), .Q(fifo_array[334])
         );
  DFFPOSX1 fifo_array_reg_20__13_ ( .D(n1048), .CLK(clk), .Q(fifo_array[333])
         );
  DFFPOSX1 fifo_array_reg_20__12_ ( .D(n1047), .CLK(clk), .Q(fifo_array[332])
         );
  DFFPOSX1 fifo_array_reg_20__11_ ( .D(n1046), .CLK(clk), .Q(fifo_array[331])
         );
  DFFPOSX1 fifo_array_reg_20__10_ ( .D(n1045), .CLK(clk), .Q(fifo_array[330])
         );
  DFFPOSX1 fifo_array_reg_20__9_ ( .D(n1044), .CLK(clk), .Q(fifo_array[329])
         );
  DFFPOSX1 fifo_array_reg_20__8_ ( .D(n1043), .CLK(clk), .Q(fifo_array[328])
         );
  DFFPOSX1 fifo_array_reg_20__7_ ( .D(n1042), .CLK(clk), .Q(fifo_array[327])
         );
  DFFPOSX1 fifo_array_reg_20__6_ ( .D(n1041), .CLK(clk), .Q(fifo_array[326])
         );
  DFFPOSX1 fifo_array_reg_20__5_ ( .D(n1040), .CLK(clk), .Q(fifo_array[325])
         );
  DFFPOSX1 fifo_array_reg_20__4_ ( .D(n1039), .CLK(clk), .Q(fifo_array[324])
         );
  DFFPOSX1 fifo_array_reg_20__3_ ( .D(n1038), .CLK(clk), .Q(fifo_array[323])
         );
  DFFPOSX1 fifo_array_reg_20__2_ ( .D(n1037), .CLK(clk), .Q(fifo_array[322])
         );
  DFFPOSX1 fifo_array_reg_20__1_ ( .D(n1036), .CLK(clk), .Q(fifo_array[321])
         );
  DFFPOSX1 fifo_array_reg_20__0_ ( .D(n1035), .CLK(clk), .Q(fifo_array[320])
         );
  DFFPOSX1 fifo_array_reg_19__15_ ( .D(n1034), .CLK(clk), .Q(fifo_array[319])
         );
  DFFPOSX1 fifo_array_reg_19__14_ ( .D(n1033), .CLK(clk), .Q(fifo_array[318])
         );
  DFFPOSX1 fifo_array_reg_19__13_ ( .D(n1032), .CLK(clk), .Q(fifo_array[317])
         );
  DFFPOSX1 fifo_array_reg_19__12_ ( .D(n1031), .CLK(clk), .Q(fifo_array[316])
         );
  DFFPOSX1 fifo_array_reg_19__11_ ( .D(n1030), .CLK(clk), .Q(fifo_array[315])
         );
  DFFPOSX1 fifo_array_reg_19__10_ ( .D(n1029), .CLK(clk), .Q(fifo_array[314])
         );
  DFFPOSX1 fifo_array_reg_19__9_ ( .D(n1028), .CLK(clk), .Q(fifo_array[313])
         );
  DFFPOSX1 fifo_array_reg_19__8_ ( .D(n1027), .CLK(clk), .Q(fifo_array[312])
         );
  DFFPOSX1 fifo_array_reg_19__7_ ( .D(n1026), .CLK(clk), .Q(fifo_array[311])
         );
  DFFPOSX1 fifo_array_reg_19__6_ ( .D(n1025), .CLK(clk), .Q(fifo_array[310])
         );
  DFFPOSX1 fifo_array_reg_19__5_ ( .D(n1024), .CLK(clk), .Q(fifo_array[309])
         );
  DFFPOSX1 fifo_array_reg_19__4_ ( .D(n1023), .CLK(clk), .Q(fifo_array[308])
         );
  DFFPOSX1 fifo_array_reg_19__3_ ( .D(n1022), .CLK(clk), .Q(fifo_array[307])
         );
  DFFPOSX1 fifo_array_reg_19__2_ ( .D(n1021), .CLK(clk), .Q(fifo_array[306])
         );
  DFFPOSX1 fifo_array_reg_19__1_ ( .D(n1020), .CLK(clk), .Q(fifo_array[305])
         );
  DFFPOSX1 fifo_array_reg_19__0_ ( .D(n1019), .CLK(clk), .Q(fifo_array[304])
         );
  DFFPOSX1 fifo_array_reg_18__15_ ( .D(n1018), .CLK(clk), .Q(fifo_array[303])
         );
  DFFPOSX1 fifo_array_reg_18__14_ ( .D(n1017), .CLK(clk), .Q(fifo_array[302])
         );
  DFFPOSX1 fifo_array_reg_18__13_ ( .D(n1016), .CLK(clk), .Q(fifo_array[301])
         );
  DFFPOSX1 fifo_array_reg_18__12_ ( .D(n1015), .CLK(clk), .Q(fifo_array[300])
         );
  DFFPOSX1 fifo_array_reg_18__11_ ( .D(n1014), .CLK(clk), .Q(fifo_array[299])
         );
  DFFPOSX1 fifo_array_reg_18__10_ ( .D(n1013), .CLK(clk), .Q(fifo_array[298])
         );
  DFFPOSX1 fifo_array_reg_18__9_ ( .D(n1012), .CLK(clk), .Q(fifo_array[297])
         );
  DFFPOSX1 fifo_array_reg_18__8_ ( .D(n1011), .CLK(clk), .Q(fifo_array[296])
         );
  DFFPOSX1 fifo_array_reg_18__7_ ( .D(n1010), .CLK(clk), .Q(fifo_array[295])
         );
  DFFPOSX1 fifo_array_reg_18__6_ ( .D(n1009), .CLK(clk), .Q(fifo_array[294])
         );
  DFFPOSX1 fifo_array_reg_18__5_ ( .D(n1008), .CLK(clk), .Q(fifo_array[293])
         );
  DFFPOSX1 fifo_array_reg_18__4_ ( .D(n1007), .CLK(clk), .Q(fifo_array[292])
         );
  DFFPOSX1 fifo_array_reg_18__3_ ( .D(n1006), .CLK(clk), .Q(fifo_array[291])
         );
  DFFPOSX1 fifo_array_reg_18__2_ ( .D(n1005), .CLK(clk), .Q(fifo_array[290])
         );
  DFFPOSX1 fifo_array_reg_18__1_ ( .D(n1004), .CLK(clk), .Q(fifo_array[289])
         );
  DFFPOSX1 fifo_array_reg_18__0_ ( .D(n1003), .CLK(clk), .Q(fifo_array[288])
         );
  DFFPOSX1 fifo_array_reg_17__15_ ( .D(n1002), .CLK(clk), .Q(fifo_array[287])
         );
  DFFPOSX1 fifo_array_reg_17__14_ ( .D(n1001), .CLK(clk), .Q(fifo_array[286])
         );
  DFFPOSX1 fifo_array_reg_17__13_ ( .D(n1000), .CLK(clk), .Q(fifo_array[285])
         );
  DFFPOSX1 fifo_array_reg_17__12_ ( .D(n999), .CLK(clk), .Q(fifo_array[284])
         );
  DFFPOSX1 fifo_array_reg_17__11_ ( .D(n998), .CLK(clk), .Q(fifo_array[283])
         );
  DFFPOSX1 fifo_array_reg_17__10_ ( .D(n997), .CLK(clk), .Q(fifo_array[282])
         );
  DFFPOSX1 fifo_array_reg_17__9_ ( .D(n996), .CLK(clk), .Q(fifo_array[281]) );
  DFFPOSX1 fifo_array_reg_17__8_ ( .D(n995), .CLK(clk), .Q(fifo_array[280]) );
  DFFPOSX1 fifo_array_reg_17__7_ ( .D(n994), .CLK(clk), .Q(fifo_array[279]) );
  DFFPOSX1 fifo_array_reg_17__6_ ( .D(n993), .CLK(clk), .Q(fifo_array[278]) );
  DFFPOSX1 fifo_array_reg_17__5_ ( .D(n992), .CLK(clk), .Q(fifo_array[277]) );
  DFFPOSX1 fifo_array_reg_17__4_ ( .D(n991), .CLK(clk), .Q(fifo_array[276]) );
  DFFPOSX1 fifo_array_reg_17__3_ ( .D(n990), .CLK(clk), .Q(fifo_array[275]) );
  DFFPOSX1 fifo_array_reg_17__2_ ( .D(n989), .CLK(clk), .Q(fifo_array[274]) );
  DFFPOSX1 fifo_array_reg_17__1_ ( .D(n988), .CLK(clk), .Q(fifo_array[273]) );
  DFFPOSX1 fifo_array_reg_17__0_ ( .D(n987), .CLK(clk), .Q(fifo_array[272]) );
  DFFPOSX1 fifo_array_reg_16__15_ ( .D(n986), .CLK(clk), .Q(fifo_array[271])
         );
  DFFPOSX1 fifo_array_reg_16__14_ ( .D(n985), .CLK(clk), .Q(fifo_array[270])
         );
  DFFPOSX1 fifo_array_reg_16__13_ ( .D(n984), .CLK(clk), .Q(fifo_array[269])
         );
  DFFPOSX1 fifo_array_reg_16__12_ ( .D(n983), .CLK(clk), .Q(fifo_array[268])
         );
  DFFPOSX1 fifo_array_reg_16__11_ ( .D(n982), .CLK(clk), .Q(fifo_array[267])
         );
  DFFPOSX1 fifo_array_reg_16__10_ ( .D(n981), .CLK(clk), .Q(fifo_array[266])
         );
  DFFPOSX1 fifo_array_reg_16__9_ ( .D(n980), .CLK(clk), .Q(fifo_array[265]) );
  DFFPOSX1 fifo_array_reg_16__8_ ( .D(n979), .CLK(clk), .Q(fifo_array[264]) );
  DFFPOSX1 fifo_array_reg_16__7_ ( .D(n978), .CLK(clk), .Q(fifo_array[263]) );
  DFFPOSX1 fifo_array_reg_16__6_ ( .D(n977), .CLK(clk), .Q(fifo_array[262]) );
  DFFPOSX1 fifo_array_reg_16__5_ ( .D(n976), .CLK(clk), .Q(fifo_array[261]) );
  DFFPOSX1 fifo_array_reg_16__4_ ( .D(n975), .CLK(clk), .Q(fifo_array[260]) );
  DFFPOSX1 fifo_array_reg_16__3_ ( .D(n974), .CLK(clk), .Q(fifo_array[259]) );
  DFFPOSX1 fifo_array_reg_16__2_ ( .D(n973), .CLK(clk), .Q(fifo_array[258]) );
  DFFPOSX1 fifo_array_reg_16__1_ ( .D(n972), .CLK(clk), .Q(fifo_array[257]) );
  DFFPOSX1 fifo_array_reg_16__0_ ( .D(n971), .CLK(clk), .Q(fifo_array[256]) );
  DFFPOSX1 fifo_array_reg_15__15_ ( .D(n970), .CLK(clk), .Q(fifo_array[255])
         );
  DFFPOSX1 fifo_array_reg_15__14_ ( .D(n969), .CLK(clk), .Q(fifo_array[254])
         );
  DFFPOSX1 fifo_array_reg_15__13_ ( .D(n968), .CLK(clk), .Q(fifo_array[253])
         );
  DFFPOSX1 fifo_array_reg_15__12_ ( .D(n967), .CLK(clk), .Q(fifo_array[252])
         );
  DFFPOSX1 fifo_array_reg_15__11_ ( .D(n966), .CLK(clk), .Q(fifo_array[251])
         );
  DFFPOSX1 fifo_array_reg_15__10_ ( .D(n965), .CLK(clk), .Q(fifo_array[250])
         );
  DFFPOSX1 fifo_array_reg_15__9_ ( .D(n964), .CLK(clk), .Q(fifo_array[249]) );
  DFFPOSX1 fifo_array_reg_15__8_ ( .D(n963), .CLK(clk), .Q(fifo_array[248]) );
  DFFPOSX1 fifo_array_reg_15__7_ ( .D(n962), .CLK(clk), .Q(fifo_array[247]) );
  DFFPOSX1 fifo_array_reg_15__6_ ( .D(n961), .CLK(clk), .Q(fifo_array[246]) );
  DFFPOSX1 fifo_array_reg_15__5_ ( .D(n960), .CLK(clk), .Q(fifo_array[245]) );
  DFFPOSX1 fifo_array_reg_15__4_ ( .D(n959), .CLK(clk), .Q(fifo_array[244]) );
  DFFPOSX1 fifo_array_reg_15__3_ ( .D(n958), .CLK(clk), .Q(fifo_array[243]) );
  DFFPOSX1 fifo_array_reg_15__2_ ( .D(n957), .CLK(clk), .Q(fifo_array[242]) );
  DFFPOSX1 fifo_array_reg_15__1_ ( .D(n956), .CLK(clk), .Q(fifo_array[241]) );
  DFFPOSX1 fifo_array_reg_15__0_ ( .D(n955), .CLK(clk), .Q(fifo_array[240]) );
  DFFPOSX1 fifo_array_reg_14__15_ ( .D(n954), .CLK(clk), .Q(fifo_array[239])
         );
  DFFPOSX1 fifo_array_reg_14__14_ ( .D(n953), .CLK(clk), .Q(fifo_array[238])
         );
  DFFPOSX1 fifo_array_reg_14__13_ ( .D(n952), .CLK(clk), .Q(fifo_array[237])
         );
  DFFPOSX1 fifo_array_reg_14__12_ ( .D(n951), .CLK(clk), .Q(fifo_array[236])
         );
  DFFPOSX1 fifo_array_reg_14__11_ ( .D(n950), .CLK(clk), .Q(fifo_array[235])
         );
  DFFPOSX1 fifo_array_reg_14__10_ ( .D(n949), .CLK(clk), .Q(fifo_array[234])
         );
  DFFPOSX1 fifo_array_reg_14__9_ ( .D(n948), .CLK(clk), .Q(fifo_array[233]) );
  DFFPOSX1 fifo_array_reg_14__8_ ( .D(n947), .CLK(clk), .Q(fifo_array[232]) );
  DFFPOSX1 fifo_array_reg_14__7_ ( .D(n946), .CLK(clk), .Q(fifo_array[231]) );
  DFFPOSX1 fifo_array_reg_14__6_ ( .D(n945), .CLK(clk), .Q(fifo_array[230]) );
  DFFPOSX1 fifo_array_reg_14__5_ ( .D(n944), .CLK(clk), .Q(fifo_array[229]) );
  DFFPOSX1 fifo_array_reg_14__4_ ( .D(n943), .CLK(clk), .Q(fifo_array[228]) );
  DFFPOSX1 fifo_array_reg_14__3_ ( .D(n942), .CLK(clk), .Q(fifo_array[227]) );
  DFFPOSX1 fifo_array_reg_14__2_ ( .D(n941), .CLK(clk), .Q(fifo_array[226]) );
  DFFPOSX1 fifo_array_reg_14__1_ ( .D(n940), .CLK(clk), .Q(fifo_array[225]) );
  DFFPOSX1 fifo_array_reg_14__0_ ( .D(n939), .CLK(clk), .Q(fifo_array[224]) );
  DFFPOSX1 fifo_array_reg_13__15_ ( .D(n938), .CLK(clk), .Q(fifo_array[223])
         );
  DFFPOSX1 fifo_array_reg_13__14_ ( .D(n937), .CLK(clk), .Q(fifo_array[222])
         );
  DFFPOSX1 fifo_array_reg_13__13_ ( .D(n936), .CLK(clk), .Q(fifo_array[221])
         );
  DFFPOSX1 fifo_array_reg_13__12_ ( .D(n935), .CLK(clk), .Q(fifo_array[220])
         );
  DFFPOSX1 fifo_array_reg_13__11_ ( .D(n934), .CLK(clk), .Q(fifo_array[219])
         );
  DFFPOSX1 fifo_array_reg_13__10_ ( .D(n933), .CLK(clk), .Q(fifo_array[218])
         );
  DFFPOSX1 fifo_array_reg_13__9_ ( .D(n932), .CLK(clk), .Q(fifo_array[217]) );
  DFFPOSX1 fifo_array_reg_13__8_ ( .D(n931), .CLK(clk), .Q(fifo_array[216]) );
  DFFPOSX1 fifo_array_reg_13__7_ ( .D(n930), .CLK(clk), .Q(fifo_array[215]) );
  DFFPOSX1 fifo_array_reg_13__6_ ( .D(n929), .CLK(clk), .Q(fifo_array[214]) );
  DFFPOSX1 fifo_array_reg_13__5_ ( .D(n928), .CLK(clk), .Q(fifo_array[213]) );
  DFFPOSX1 fifo_array_reg_13__4_ ( .D(n927), .CLK(clk), .Q(fifo_array[212]) );
  DFFPOSX1 fifo_array_reg_13__3_ ( .D(n926), .CLK(clk), .Q(fifo_array[211]) );
  DFFPOSX1 fifo_array_reg_13__2_ ( .D(n925), .CLK(clk), .Q(fifo_array[210]) );
  DFFPOSX1 fifo_array_reg_13__1_ ( .D(n924), .CLK(clk), .Q(fifo_array[209]) );
  DFFPOSX1 fifo_array_reg_13__0_ ( .D(n923), .CLK(clk), .Q(fifo_array[208]) );
  DFFPOSX1 fifo_array_reg_12__15_ ( .D(n922), .CLK(clk), .Q(fifo_array[207])
         );
  DFFPOSX1 fifo_array_reg_12__14_ ( .D(n921), .CLK(clk), .Q(fifo_array[206])
         );
  DFFPOSX1 fifo_array_reg_12__13_ ( .D(n920), .CLK(clk), .Q(fifo_array[205])
         );
  DFFPOSX1 fifo_array_reg_12__12_ ( .D(n919), .CLK(clk), .Q(fifo_array[204])
         );
  DFFPOSX1 fifo_array_reg_12__11_ ( .D(n918), .CLK(clk), .Q(fifo_array[203])
         );
  DFFPOSX1 fifo_array_reg_12__10_ ( .D(n917), .CLK(clk), .Q(fifo_array[202])
         );
  DFFPOSX1 fifo_array_reg_12__9_ ( .D(n916), .CLK(clk), .Q(fifo_array[201]) );
  DFFPOSX1 fifo_array_reg_12__8_ ( .D(n915), .CLK(clk), .Q(fifo_array[200]) );
  DFFPOSX1 fifo_array_reg_12__7_ ( .D(n914), .CLK(clk), .Q(fifo_array[199]) );
  DFFPOSX1 fifo_array_reg_12__6_ ( .D(n913), .CLK(clk), .Q(fifo_array[198]) );
  DFFPOSX1 fifo_array_reg_12__5_ ( .D(n912), .CLK(clk), .Q(fifo_array[197]) );
  DFFPOSX1 fifo_array_reg_12__4_ ( .D(n911), .CLK(clk), .Q(fifo_array[196]) );
  DFFPOSX1 fifo_array_reg_12__3_ ( .D(n910), .CLK(clk), .Q(fifo_array[195]) );
  DFFPOSX1 fifo_array_reg_12__2_ ( .D(n909), .CLK(clk), .Q(fifo_array[194]) );
  DFFPOSX1 fifo_array_reg_12__1_ ( .D(n908), .CLK(clk), .Q(fifo_array[193]) );
  DFFPOSX1 fifo_array_reg_12__0_ ( .D(n907), .CLK(clk), .Q(fifo_array[192]) );
  DFFPOSX1 fifo_array_reg_11__15_ ( .D(n906), .CLK(clk), .Q(fifo_array[191])
         );
  DFFPOSX1 fifo_array_reg_11__14_ ( .D(n905), .CLK(clk), .Q(fifo_array[190])
         );
  DFFPOSX1 fifo_array_reg_11__13_ ( .D(n904), .CLK(clk), .Q(fifo_array[189])
         );
  DFFPOSX1 fifo_array_reg_11__12_ ( .D(n903), .CLK(clk), .Q(fifo_array[188])
         );
  DFFPOSX1 fifo_array_reg_11__11_ ( .D(n902), .CLK(clk), .Q(fifo_array[187])
         );
  DFFPOSX1 fifo_array_reg_11__10_ ( .D(n901), .CLK(clk), .Q(fifo_array[186])
         );
  DFFPOSX1 fifo_array_reg_11__9_ ( .D(n900), .CLK(clk), .Q(fifo_array[185]) );
  DFFPOSX1 fifo_array_reg_11__8_ ( .D(n899), .CLK(clk), .Q(fifo_array[184]) );
  DFFPOSX1 fifo_array_reg_11__7_ ( .D(n898), .CLK(clk), .Q(fifo_array[183]) );
  DFFPOSX1 fifo_array_reg_11__6_ ( .D(n897), .CLK(clk), .Q(fifo_array[182]) );
  DFFPOSX1 fifo_array_reg_11__5_ ( .D(n896), .CLK(clk), .Q(fifo_array[181]) );
  DFFPOSX1 fifo_array_reg_11__4_ ( .D(n895), .CLK(clk), .Q(fifo_array[180]) );
  DFFPOSX1 fifo_array_reg_11__3_ ( .D(n894), .CLK(clk), .Q(fifo_array[179]) );
  DFFPOSX1 fifo_array_reg_11__2_ ( .D(n893), .CLK(clk), .Q(fifo_array[178]) );
  DFFPOSX1 fifo_array_reg_11__1_ ( .D(n892), .CLK(clk), .Q(fifo_array[177]) );
  DFFPOSX1 fifo_array_reg_11__0_ ( .D(n891), .CLK(clk), .Q(fifo_array[176]) );
  DFFPOSX1 fifo_array_reg_10__15_ ( .D(n890), .CLK(clk), .Q(fifo_array[175])
         );
  DFFPOSX1 fifo_array_reg_10__14_ ( .D(n889), .CLK(clk), .Q(fifo_array[174])
         );
  DFFPOSX1 fifo_array_reg_10__13_ ( .D(n888), .CLK(clk), .Q(fifo_array[173])
         );
  DFFPOSX1 fifo_array_reg_10__12_ ( .D(n887), .CLK(clk), .Q(fifo_array[172])
         );
  DFFPOSX1 fifo_array_reg_10__11_ ( .D(n886), .CLK(clk), .Q(fifo_array[171])
         );
  DFFPOSX1 fifo_array_reg_10__10_ ( .D(n885), .CLK(clk), .Q(fifo_array[170])
         );
  DFFPOSX1 fifo_array_reg_10__9_ ( .D(n884), .CLK(clk), .Q(fifo_array[169]) );
  DFFPOSX1 fifo_array_reg_10__8_ ( .D(n883), .CLK(clk), .Q(fifo_array[168]) );
  DFFPOSX1 fifo_array_reg_10__7_ ( .D(n882), .CLK(clk), .Q(fifo_array[167]) );
  DFFPOSX1 fifo_array_reg_10__6_ ( .D(n881), .CLK(clk), .Q(fifo_array[166]) );
  DFFPOSX1 fifo_array_reg_10__5_ ( .D(n880), .CLK(clk), .Q(fifo_array[165]) );
  DFFPOSX1 fifo_array_reg_10__4_ ( .D(n879), .CLK(clk), .Q(fifo_array[164]) );
  DFFPOSX1 fifo_array_reg_10__3_ ( .D(n878), .CLK(clk), .Q(fifo_array[163]) );
  DFFPOSX1 fifo_array_reg_10__2_ ( .D(n877), .CLK(clk), .Q(fifo_array[162]) );
  DFFPOSX1 fifo_array_reg_10__1_ ( .D(n876), .CLK(clk), .Q(fifo_array[161]) );
  DFFPOSX1 fifo_array_reg_10__0_ ( .D(n875), .CLK(clk), .Q(fifo_array[160]) );
  DFFPOSX1 fifo_array_reg_9__15_ ( .D(n874), .CLK(clk), .Q(fifo_array[159]) );
  DFFPOSX1 fifo_array_reg_9__14_ ( .D(n873), .CLK(clk), .Q(fifo_array[158]) );
  DFFPOSX1 fifo_array_reg_9__13_ ( .D(n872), .CLK(clk), .Q(fifo_array[157]) );
  DFFPOSX1 fifo_array_reg_9__12_ ( .D(n871), .CLK(clk), .Q(fifo_array[156]) );
  DFFPOSX1 fifo_array_reg_9__11_ ( .D(n870), .CLK(clk), .Q(fifo_array[155]) );
  DFFPOSX1 fifo_array_reg_9__10_ ( .D(n869), .CLK(clk), .Q(fifo_array[154]) );
  DFFPOSX1 fifo_array_reg_9__9_ ( .D(n868), .CLK(clk), .Q(fifo_array[153]) );
  DFFPOSX1 fifo_array_reg_9__8_ ( .D(n867), .CLK(clk), .Q(fifo_array[152]) );
  DFFPOSX1 fifo_array_reg_9__7_ ( .D(n866), .CLK(clk), .Q(fifo_array[151]) );
  DFFPOSX1 fifo_array_reg_9__6_ ( .D(n865), .CLK(clk), .Q(fifo_array[150]) );
  DFFPOSX1 fifo_array_reg_9__5_ ( .D(n864), .CLK(clk), .Q(fifo_array[149]) );
  DFFPOSX1 fifo_array_reg_9__4_ ( .D(n863), .CLK(clk), .Q(fifo_array[148]) );
  DFFPOSX1 fifo_array_reg_9__3_ ( .D(n862), .CLK(clk), .Q(fifo_array[147]) );
  DFFPOSX1 fifo_array_reg_9__2_ ( .D(n861), .CLK(clk), .Q(fifo_array[146]) );
  DFFPOSX1 fifo_array_reg_9__1_ ( .D(n860), .CLK(clk), .Q(fifo_array[145]) );
  DFFPOSX1 fifo_array_reg_9__0_ ( .D(n859), .CLK(clk), .Q(fifo_array[144]) );
  DFFPOSX1 fifo_array_reg_8__15_ ( .D(n858), .CLK(clk), .Q(fifo_array[143]) );
  DFFPOSX1 fifo_array_reg_8__14_ ( .D(n857), .CLK(clk), .Q(fifo_array[142]) );
  DFFPOSX1 fifo_array_reg_8__13_ ( .D(n856), .CLK(clk), .Q(fifo_array[141]) );
  DFFPOSX1 fifo_array_reg_8__12_ ( .D(n855), .CLK(clk), .Q(fifo_array[140]) );
  DFFPOSX1 fifo_array_reg_8__11_ ( .D(n854), .CLK(clk), .Q(fifo_array[139]) );
  DFFPOSX1 fifo_array_reg_8__10_ ( .D(n853), .CLK(clk), .Q(fifo_array[138]) );
  DFFPOSX1 fifo_array_reg_8__9_ ( .D(n852), .CLK(clk), .Q(fifo_array[137]) );
  DFFPOSX1 fifo_array_reg_8__8_ ( .D(n851), .CLK(clk), .Q(fifo_array[136]) );
  DFFPOSX1 fifo_array_reg_8__7_ ( .D(n850), .CLK(clk), .Q(fifo_array[135]) );
  DFFPOSX1 fifo_array_reg_8__6_ ( .D(n849), .CLK(clk), .Q(fifo_array[134]) );
  DFFPOSX1 fifo_array_reg_8__5_ ( .D(n848), .CLK(clk), .Q(fifo_array[133]) );
  DFFPOSX1 fifo_array_reg_8__4_ ( .D(n847), .CLK(clk), .Q(fifo_array[132]) );
  DFFPOSX1 fifo_array_reg_8__3_ ( .D(n846), .CLK(clk), .Q(fifo_array[131]) );
  DFFPOSX1 fifo_array_reg_8__2_ ( .D(n845), .CLK(clk), .Q(fifo_array[130]) );
  DFFPOSX1 fifo_array_reg_8__1_ ( .D(n844), .CLK(clk), .Q(fifo_array[129]) );
  DFFPOSX1 fifo_array_reg_8__0_ ( .D(n843), .CLK(clk), .Q(fifo_array[128]) );
  DFFPOSX1 fifo_array_reg_7__15_ ( .D(n842), .CLK(clk), .Q(fifo_array[127]) );
  DFFPOSX1 fifo_array_reg_7__14_ ( .D(n841), .CLK(clk), .Q(fifo_array[126]) );
  DFFPOSX1 fifo_array_reg_7__13_ ( .D(n840), .CLK(clk), .Q(fifo_array[125]) );
  DFFPOSX1 fifo_array_reg_7__12_ ( .D(n839), .CLK(clk), .Q(fifo_array[124]) );
  DFFPOSX1 fifo_array_reg_7__11_ ( .D(n838), .CLK(clk), .Q(fifo_array[123]) );
  DFFPOSX1 fifo_array_reg_7__10_ ( .D(n837), .CLK(clk), .Q(fifo_array[122]) );
  DFFPOSX1 fifo_array_reg_7__9_ ( .D(n836), .CLK(clk), .Q(fifo_array[121]) );
  DFFPOSX1 fifo_array_reg_7__8_ ( .D(n835), .CLK(clk), .Q(fifo_array[120]) );
  DFFPOSX1 fifo_array_reg_7__7_ ( .D(n834), .CLK(clk), .Q(fifo_array[119]) );
  DFFPOSX1 fifo_array_reg_7__6_ ( .D(n833), .CLK(clk), .Q(fifo_array[118]) );
  DFFPOSX1 fifo_array_reg_7__5_ ( .D(n832), .CLK(clk), .Q(fifo_array[117]) );
  DFFPOSX1 fifo_array_reg_7__4_ ( .D(n831), .CLK(clk), .Q(fifo_array[116]) );
  DFFPOSX1 fifo_array_reg_7__3_ ( .D(n830), .CLK(clk), .Q(fifo_array[115]) );
  DFFPOSX1 fifo_array_reg_7__2_ ( .D(n829), .CLK(clk), .Q(fifo_array[114]) );
  DFFPOSX1 fifo_array_reg_7__1_ ( .D(n828), .CLK(clk), .Q(fifo_array[113]) );
  DFFPOSX1 fifo_array_reg_7__0_ ( .D(n827), .CLK(clk), .Q(fifo_array[112]) );
  DFFPOSX1 fifo_array_reg_6__15_ ( .D(n826), .CLK(clk), .Q(fifo_array[111]) );
  DFFPOSX1 fifo_array_reg_6__14_ ( .D(n825), .CLK(clk), .Q(fifo_array[110]) );
  DFFPOSX1 fifo_array_reg_6__13_ ( .D(n824), .CLK(clk), .Q(fifo_array[109]) );
  DFFPOSX1 fifo_array_reg_6__12_ ( .D(n823), .CLK(clk), .Q(fifo_array[108]) );
  DFFPOSX1 fifo_array_reg_6__11_ ( .D(n822), .CLK(clk), .Q(fifo_array[107]) );
  DFFPOSX1 fifo_array_reg_6__10_ ( .D(n821), .CLK(clk), .Q(fifo_array[106]) );
  DFFPOSX1 fifo_array_reg_6__9_ ( .D(n820), .CLK(clk), .Q(fifo_array[105]) );
  DFFPOSX1 fifo_array_reg_6__8_ ( .D(n819), .CLK(clk), .Q(fifo_array[104]) );
  DFFPOSX1 fifo_array_reg_6__7_ ( .D(n818), .CLK(clk), .Q(fifo_array[103]) );
  DFFPOSX1 fifo_array_reg_6__6_ ( .D(n817), .CLK(clk), .Q(fifo_array[102]) );
  DFFPOSX1 fifo_array_reg_6__5_ ( .D(n816), .CLK(clk), .Q(fifo_array[101]) );
  DFFPOSX1 fifo_array_reg_6__4_ ( .D(n815), .CLK(clk), .Q(fifo_array[100]) );
  DFFPOSX1 fifo_array_reg_6__3_ ( .D(n814), .CLK(clk), .Q(fifo_array[99]) );
  DFFPOSX1 fifo_array_reg_6__2_ ( .D(n813), .CLK(clk), .Q(fifo_array[98]) );
  DFFPOSX1 fifo_array_reg_6__1_ ( .D(n812), .CLK(clk), .Q(fifo_array[97]) );
  DFFPOSX1 fifo_array_reg_6__0_ ( .D(n811), .CLK(clk), .Q(fifo_array[96]) );
  DFFPOSX1 fifo_array_reg_5__15_ ( .D(n810), .CLK(clk), .Q(fifo_array[95]) );
  DFFPOSX1 fifo_array_reg_5__14_ ( .D(n809), .CLK(clk), .Q(fifo_array[94]) );
  DFFPOSX1 fifo_array_reg_5__13_ ( .D(n808), .CLK(clk), .Q(fifo_array[93]) );
  DFFPOSX1 fifo_array_reg_5__12_ ( .D(n807), .CLK(clk), .Q(fifo_array[92]) );
  DFFPOSX1 fifo_array_reg_5__11_ ( .D(n806), .CLK(clk), .Q(fifo_array[91]) );
  DFFPOSX1 fifo_array_reg_5__10_ ( .D(n805), .CLK(clk), .Q(fifo_array[90]) );
  DFFPOSX1 fifo_array_reg_5__9_ ( .D(n804), .CLK(clk), .Q(fifo_array[89]) );
  DFFPOSX1 fifo_array_reg_5__8_ ( .D(n803), .CLK(clk), .Q(fifo_array[88]) );
  DFFPOSX1 fifo_array_reg_5__7_ ( .D(n802), .CLK(clk), .Q(fifo_array[87]) );
  DFFPOSX1 fifo_array_reg_5__6_ ( .D(n801), .CLK(clk), .Q(fifo_array[86]) );
  DFFPOSX1 fifo_array_reg_5__5_ ( .D(n800), .CLK(clk), .Q(fifo_array[85]) );
  DFFPOSX1 fifo_array_reg_5__4_ ( .D(n799), .CLK(clk), .Q(fifo_array[84]) );
  DFFPOSX1 fifo_array_reg_5__3_ ( .D(n798), .CLK(clk), .Q(fifo_array[83]) );
  DFFPOSX1 fifo_array_reg_5__2_ ( .D(n797), .CLK(clk), .Q(fifo_array[82]) );
  DFFPOSX1 fifo_array_reg_5__1_ ( .D(n796), .CLK(clk), .Q(fifo_array[81]) );
  DFFPOSX1 fifo_array_reg_5__0_ ( .D(n795), .CLK(clk), .Q(fifo_array[80]) );
  DFFPOSX1 fifo_array_reg_4__15_ ( .D(n794), .CLK(clk), .Q(fifo_array[79]) );
  DFFPOSX1 fifo_array_reg_4__14_ ( .D(n793), .CLK(clk), .Q(fifo_array[78]) );
  DFFPOSX1 fifo_array_reg_4__13_ ( .D(n792), .CLK(clk), .Q(fifo_array[77]) );
  DFFPOSX1 fifo_array_reg_4__12_ ( .D(n791), .CLK(clk), .Q(fifo_array[76]) );
  DFFPOSX1 fifo_array_reg_4__11_ ( .D(n790), .CLK(clk), .Q(fifo_array[75]) );
  DFFPOSX1 fifo_array_reg_4__10_ ( .D(n789), .CLK(clk), .Q(fifo_array[74]) );
  DFFPOSX1 fifo_array_reg_4__9_ ( .D(n788), .CLK(clk), .Q(fifo_array[73]) );
  DFFPOSX1 fifo_array_reg_4__8_ ( .D(n787), .CLK(clk), .Q(fifo_array[72]) );
  DFFPOSX1 fifo_array_reg_4__7_ ( .D(n786), .CLK(clk), .Q(fifo_array[71]) );
  DFFPOSX1 fifo_array_reg_4__6_ ( .D(n785), .CLK(clk), .Q(fifo_array[70]) );
  DFFPOSX1 fifo_array_reg_4__5_ ( .D(n784), .CLK(clk), .Q(fifo_array[69]) );
  DFFPOSX1 fifo_array_reg_4__4_ ( .D(n783), .CLK(clk), .Q(fifo_array[68]) );
  DFFPOSX1 fifo_array_reg_4__3_ ( .D(n782), .CLK(clk), .Q(fifo_array[67]) );
  DFFPOSX1 fifo_array_reg_4__2_ ( .D(n781), .CLK(clk), .Q(fifo_array[66]) );
  DFFPOSX1 fifo_array_reg_4__1_ ( .D(n780), .CLK(clk), .Q(fifo_array[65]) );
  DFFPOSX1 fifo_array_reg_4__0_ ( .D(n779), .CLK(clk), .Q(fifo_array[64]) );
  DFFPOSX1 fifo_array_reg_3__15_ ( .D(n778), .CLK(clk), .Q(fifo_array[63]) );
  DFFPOSX1 fifo_array_reg_3__14_ ( .D(n777), .CLK(clk), .Q(fifo_array[62]) );
  DFFPOSX1 fifo_array_reg_3__13_ ( .D(n776), .CLK(clk), .Q(fifo_array[61]) );
  DFFPOSX1 fifo_array_reg_3__12_ ( .D(n775), .CLK(clk), .Q(fifo_array[60]) );
  DFFPOSX1 fifo_array_reg_3__11_ ( .D(n774), .CLK(clk), .Q(fifo_array[59]) );
  DFFPOSX1 fifo_array_reg_3__10_ ( .D(n773), .CLK(clk), .Q(fifo_array[58]) );
  DFFPOSX1 fifo_array_reg_3__9_ ( .D(n772), .CLK(clk), .Q(fifo_array[57]) );
  DFFPOSX1 fifo_array_reg_3__8_ ( .D(n771), .CLK(clk), .Q(fifo_array[56]) );
  DFFPOSX1 fifo_array_reg_3__7_ ( .D(n770), .CLK(clk), .Q(fifo_array[55]) );
  DFFPOSX1 fifo_array_reg_3__6_ ( .D(n769), .CLK(clk), .Q(fifo_array[54]) );
  DFFPOSX1 fifo_array_reg_3__5_ ( .D(n768), .CLK(clk), .Q(fifo_array[53]) );
  DFFPOSX1 fifo_array_reg_3__4_ ( .D(n767), .CLK(clk), .Q(fifo_array[52]) );
  DFFPOSX1 fifo_array_reg_3__3_ ( .D(n766), .CLK(clk), .Q(fifo_array[51]) );
  DFFPOSX1 fifo_array_reg_3__2_ ( .D(n765), .CLK(clk), .Q(fifo_array[50]) );
  DFFPOSX1 fifo_array_reg_3__1_ ( .D(n764), .CLK(clk), .Q(fifo_array[49]) );
  DFFPOSX1 fifo_array_reg_3__0_ ( .D(n763), .CLK(clk), .Q(fifo_array[48]) );
  DFFPOSX1 fifo_array_reg_2__15_ ( .D(n762), .CLK(clk), .Q(fifo_array[47]) );
  DFFPOSX1 fifo_array_reg_2__14_ ( .D(n761), .CLK(clk), .Q(fifo_array[46]) );
  DFFPOSX1 fifo_array_reg_2__13_ ( .D(n760), .CLK(clk), .Q(fifo_array[45]) );
  DFFPOSX1 fifo_array_reg_2__12_ ( .D(n759), .CLK(clk), .Q(fifo_array[44]) );
  DFFPOSX1 fifo_array_reg_2__11_ ( .D(n758), .CLK(clk), .Q(fifo_array[43]) );
  DFFPOSX1 fifo_array_reg_2__10_ ( .D(n757), .CLK(clk), .Q(fifo_array[42]) );
  DFFPOSX1 fifo_array_reg_2__9_ ( .D(n756), .CLK(clk), .Q(fifo_array[41]) );
  DFFPOSX1 fifo_array_reg_2__8_ ( .D(n755), .CLK(clk), .Q(fifo_array[40]) );
  DFFPOSX1 fifo_array_reg_2__7_ ( .D(n754), .CLK(clk), .Q(fifo_array[39]) );
  DFFPOSX1 fifo_array_reg_2__6_ ( .D(n753), .CLK(clk), .Q(fifo_array[38]) );
  DFFPOSX1 fifo_array_reg_2__5_ ( .D(n752), .CLK(clk), .Q(fifo_array[37]) );
  DFFPOSX1 fifo_array_reg_2__4_ ( .D(n751), .CLK(clk), .Q(fifo_array[36]) );
  DFFPOSX1 fifo_array_reg_2__3_ ( .D(n750), .CLK(clk), .Q(fifo_array[35]) );
  DFFPOSX1 fifo_array_reg_2__2_ ( .D(n749), .CLK(clk), .Q(fifo_array[34]) );
  DFFPOSX1 fifo_array_reg_2__1_ ( .D(n748), .CLK(clk), .Q(fifo_array[33]) );
  DFFPOSX1 fifo_array_reg_2__0_ ( .D(n747), .CLK(clk), .Q(fifo_array[32]) );
  DFFPOSX1 fifo_array_reg_1__15_ ( .D(n746), .CLK(clk), .Q(fifo_array[31]) );
  DFFPOSX1 fifo_array_reg_1__14_ ( .D(n745), .CLK(clk), .Q(fifo_array[30]) );
  DFFPOSX1 fifo_array_reg_1__13_ ( .D(n744), .CLK(clk), .Q(fifo_array[29]) );
  DFFPOSX1 fifo_array_reg_1__12_ ( .D(n743), .CLK(clk), .Q(fifo_array[28]) );
  DFFPOSX1 fifo_array_reg_1__11_ ( .D(n742), .CLK(clk), .Q(fifo_array[27]) );
  DFFPOSX1 fifo_array_reg_1__10_ ( .D(n741), .CLK(clk), .Q(fifo_array[26]) );
  DFFPOSX1 fifo_array_reg_1__9_ ( .D(n740), .CLK(clk), .Q(fifo_array[25]) );
  DFFPOSX1 fifo_array_reg_1__8_ ( .D(n739), .CLK(clk), .Q(fifo_array[24]) );
  DFFPOSX1 fifo_array_reg_1__7_ ( .D(n738), .CLK(clk), .Q(fifo_array[23]) );
  DFFPOSX1 fifo_array_reg_1__6_ ( .D(n737), .CLK(clk), .Q(fifo_array[22]) );
  DFFPOSX1 fifo_array_reg_1__5_ ( .D(n736), .CLK(clk), .Q(fifo_array[21]) );
  DFFPOSX1 fifo_array_reg_1__4_ ( .D(n735), .CLK(clk), .Q(fifo_array[20]) );
  DFFPOSX1 fifo_array_reg_1__3_ ( .D(n734), .CLK(clk), .Q(fifo_array[19]) );
  DFFPOSX1 fifo_array_reg_1__2_ ( .D(n733), .CLK(clk), .Q(fifo_array[18]) );
  DFFPOSX1 fifo_array_reg_1__1_ ( .D(n732), .CLK(clk), .Q(fifo_array[17]) );
  DFFPOSX1 fifo_array_reg_1__0_ ( .D(n731), .CLK(clk), .Q(fifo_array[16]) );
  DFFPOSX1 fifo_array_reg_0__15_ ( .D(n730), .CLK(clk), .Q(fifo_array[15]) );
  DFFPOSX1 fifo_array_reg_0__14_ ( .D(n729), .CLK(clk), .Q(fifo_array[14]) );
  DFFPOSX1 fifo_array_reg_0__13_ ( .D(n728), .CLK(clk), .Q(fifo_array[13]) );
  DFFPOSX1 fifo_array_reg_0__12_ ( .D(n727), .CLK(clk), .Q(fifo_array[12]) );
  DFFPOSX1 fifo_array_reg_0__11_ ( .D(n726), .CLK(clk), .Q(fifo_array[11]) );
  DFFPOSX1 fifo_array_reg_0__10_ ( .D(n725), .CLK(clk), .Q(fifo_array[10]) );
  DFFPOSX1 fifo_array_reg_0__9_ ( .D(n724), .CLK(clk), .Q(fifo_array[9]) );
  DFFPOSX1 fifo_array_reg_0__8_ ( .D(n723), .CLK(clk), .Q(fifo_array[8]) );
  DFFPOSX1 fifo_array_reg_0__7_ ( .D(n722), .CLK(clk), .Q(fifo_array[7]) );
  DFFPOSX1 fifo_array_reg_0__6_ ( .D(n721), .CLK(clk), .Q(fifo_array[6]) );
  DFFPOSX1 fifo_array_reg_0__5_ ( .D(n720), .CLK(clk), .Q(fifo_array[5]) );
  DFFPOSX1 fifo_array_reg_0__4_ ( .D(n719), .CLK(clk), .Q(fifo_array[4]) );
  DFFPOSX1 fifo_array_reg_0__3_ ( .D(n718), .CLK(clk), .Q(fifo_array[3]) );
  DFFPOSX1 fifo_array_reg_0__2_ ( .D(n717), .CLK(clk), .Q(fifo_array[2]) );
  DFFPOSX1 fifo_array_reg_0__1_ ( .D(n716), .CLK(clk), .Q(fifo_array[1]) );
  DFFPOSX1 fifo_array_reg_0__0_ ( .D(n715), .CLK(clk), .Q(fifo_array[0]) );
  OAI21X1 U67 ( .A(n2310), .B(n2278), .C(n1706), .Y(n715) );
  OAI21X1 U69 ( .A(n2310), .B(n2277), .C(n1663), .Y(n716) );
  OAI21X1 U71 ( .A(n2310), .B(n2276), .C(n1622), .Y(n717) );
  OAI21X1 U73 ( .A(n2310), .B(n2275), .C(n1581), .Y(n718) );
  OAI21X1 U75 ( .A(n2310), .B(n2274), .C(n1539), .Y(n719) );
  OAI21X1 U77 ( .A(n2310), .B(n2273), .C(n1503), .Y(n720) );
  OAI21X1 U79 ( .A(n2310), .B(n2272), .C(n1468), .Y(n721) );
  OAI21X1 U81 ( .A(n2310), .B(n2271), .C(n1434), .Y(n722) );
  OAI21X1 U83 ( .A(n2310), .B(n2270), .C(n1400), .Y(n723) );
  OAI21X1 U85 ( .A(n2310), .B(n2269), .C(n1368), .Y(n724) );
  OAI21X1 U87 ( .A(n2310), .B(n2268), .C(n1336), .Y(n725) );
  OAI21X1 U89 ( .A(n2310), .B(n2267), .C(n1306), .Y(n726) );
  OAI21X1 U91 ( .A(n2310), .B(n2266), .C(n1705), .Y(n727) );
  OAI21X1 U93 ( .A(n2310), .B(n2265), .C(n1662), .Y(n728) );
  OAI21X1 U95 ( .A(n2310), .B(n2264), .C(n1276), .Y(n729) );
  OAI21X1 U97 ( .A(n2310), .B(n2263), .C(n1248), .Y(n730) );
  OAI21X1 U100 ( .A(n2278), .B(n2309), .C(n1661), .Y(n731) );
  OAI21X1 U102 ( .A(n2277), .B(n2309), .C(n1704), .Y(n732) );
  OAI21X1 U104 ( .A(n2276), .B(n2309), .C(n1580), .Y(n733) );
  OAI21X1 U106 ( .A(n2275), .B(n2309), .C(n1621), .Y(n734) );
  OAI21X1 U108 ( .A(n2274), .B(n2309), .C(n1502), .Y(n735) );
  OAI21X1 U110 ( .A(n2273), .B(n2309), .C(n1538), .Y(n736) );
  OAI21X1 U112 ( .A(n2272), .B(n2309), .C(n1433), .Y(n737) );
  OAI21X1 U114 ( .A(n2271), .B(n2309), .C(n1467), .Y(n738) );
  OAI21X1 U116 ( .A(n2270), .B(n2309), .C(n1367), .Y(n739) );
  OAI21X1 U118 ( .A(n2269), .B(n2309), .C(n1399), .Y(n740) );
  OAI21X1 U120 ( .A(n2268), .B(n2309), .C(n1305), .Y(n741) );
  OAI21X1 U122 ( .A(n2267), .B(n2309), .C(n1335), .Y(n742) );
  OAI21X1 U124 ( .A(n2266), .B(n2309), .C(n1660), .Y(n743) );
  OAI21X1 U126 ( .A(n2265), .B(n2309), .C(n1703), .Y(n744) );
  OAI21X1 U128 ( .A(n2264), .B(n2309), .C(n1247), .Y(n745) );
  OAI21X1 U130 ( .A(n2263), .B(n2309), .C(n1275), .Y(n746) );
  OAI21X1 U133 ( .A(n2278), .B(n2308), .C(n1620), .Y(n747) );
  OAI21X1 U135 ( .A(n2277), .B(n2308), .C(n1579), .Y(n748) );
  OAI21X1 U137 ( .A(n2276), .B(n2308), .C(n1702), .Y(n749) );
  OAI21X1 U139 ( .A(n2275), .B(n2308), .C(n1659), .Y(n750) );
  OAI21X1 U141 ( .A(n2274), .B(n2308), .C(n1466), .Y(n751) );
  OAI21X1 U143 ( .A(n2273), .B(n2308), .C(n1432), .Y(n752) );
  OAI21X1 U145 ( .A(n2272), .B(n2308), .C(n1537), .Y(n753) );
  OAI21X1 U147 ( .A(n2271), .B(n2308), .C(n1501), .Y(n754) );
  OAI21X1 U149 ( .A(n2270), .B(n2308), .C(n1334), .Y(n755) );
  OAI21X1 U151 ( .A(n2269), .B(n2308), .C(n1304), .Y(n756) );
  OAI21X1 U153 ( .A(n2268), .B(n2308), .C(n1398), .Y(n757) );
  OAI21X1 U155 ( .A(n2267), .B(n2308), .C(n1366), .Y(n758) );
  OAI21X1 U157 ( .A(n2266), .B(n2308), .C(n1619), .Y(n759) );
  OAI21X1 U159 ( .A(n2265), .B(n2308), .C(n1578), .Y(n760) );
  OAI21X1 U161 ( .A(n2264), .B(n2308), .C(n331), .Y(n761) );
  OAI21X1 U163 ( .A(n2263), .B(n2308), .C(n87), .Y(n762) );
  OAI21X1 U166 ( .A(n2278), .B(n2307), .C(n1577), .Y(n763) );
  OAI21X1 U168 ( .A(n2277), .B(n2307), .C(n1618), .Y(n764) );
  OAI21X1 U170 ( .A(n2276), .B(n2307), .C(n1658), .Y(n765) );
  OAI21X1 U172 ( .A(n2275), .B(n2307), .C(n1701), .Y(n766) );
  OAI21X1 U174 ( .A(n2274), .B(n2307), .C(n1431), .Y(n767) );
  OAI21X1 U176 ( .A(n2273), .B(n2307), .C(n1465), .Y(n768) );
  OAI21X1 U178 ( .A(n2272), .B(n2307), .C(n1500), .Y(n769) );
  OAI21X1 U180 ( .A(n2271), .B(n2307), .C(n1536), .Y(n770) );
  OAI21X1 U182 ( .A(n2270), .B(n2307), .C(n1303), .Y(n771) );
  OAI21X1 U184 ( .A(n2269), .B(n2307), .C(n1333), .Y(n772) );
  OAI21X1 U186 ( .A(n2268), .B(n2307), .C(n1365), .Y(n773) );
  OAI21X1 U188 ( .A(n2267), .B(n2307), .C(n1397), .Y(n774) );
  OAI21X1 U190 ( .A(n2266), .B(n2307), .C(n1576), .Y(n775) );
  OAI21X1 U192 ( .A(n2265), .B(n2307), .C(n1617), .Y(n776) );
  OAI21X1 U194 ( .A(n2264), .B(n2307), .C(n86), .Y(n777) );
  OAI21X1 U196 ( .A(n2263), .B(n2307), .C(n314), .Y(n778) );
  OAI21X1 U199 ( .A(n2278), .B(n2306), .C(n1535), .Y(n779) );
  OAI21X1 U201 ( .A(n2277), .B(n2306), .C(n1499), .Y(n780) );
  OAI21X1 U203 ( .A(n2276), .B(n2306), .C(n1464), .Y(n781) );
  OAI21X1 U205 ( .A(n2275), .B(n2306), .C(n1430), .Y(n782) );
  OAI21X1 U207 ( .A(n2274), .B(n2306), .C(n1700), .Y(n783) );
  OAI21X1 U209 ( .A(n2273), .B(n2306), .C(n1657), .Y(n784) );
  OAI21X1 U211 ( .A(n2272), .B(n2306), .C(n1616), .Y(n785) );
  OAI21X1 U213 ( .A(n2271), .B(n2306), .C(n1575), .Y(n786) );
  OAI21X1 U215 ( .A(n2270), .B(n2306), .C(n1274), .Y(n787) );
  OAI21X1 U217 ( .A(n2269), .B(n2306), .C(n1246), .Y(n788) );
  OAI21X1 U219 ( .A(n2268), .B(n2306), .C(n297), .Y(n789) );
  OAI21X1 U221 ( .A(n2267), .B(n2306), .C(n85), .Y(n790) );
  OAI21X1 U223 ( .A(n2266), .B(n2306), .C(n1534), .Y(n791) );
  OAI21X1 U225 ( .A(n2265), .B(n2306), .C(n1498), .Y(n792) );
  OAI21X1 U227 ( .A(n2264), .B(n2306), .C(n1396), .Y(n793) );
  OAI21X1 U229 ( .A(n2263), .B(n2306), .C(n1364), .Y(n794) );
  OAI21X1 U232 ( .A(n2278), .B(n2305), .C(n1497), .Y(n795) );
  OAI21X1 U234 ( .A(n2277), .B(n2305), .C(n1533), .Y(n796) );
  OAI21X1 U236 ( .A(n2276), .B(n2305), .C(n1429), .Y(n797) );
  OAI21X1 U238 ( .A(n2275), .B(n2305), .C(n1463), .Y(n798) );
  OAI21X1 U240 ( .A(n2274), .B(n2305), .C(n1656), .Y(n799) );
  OAI21X1 U242 ( .A(n2273), .B(n2305), .C(n1699), .Y(n800) );
  OAI21X1 U244 ( .A(n2272), .B(n2305), .C(n1574), .Y(n801) );
  OAI21X1 U246 ( .A(n2271), .B(n2305), .C(n1615), .Y(n802) );
  OAI21X1 U248 ( .A(n2270), .B(n2305), .C(n1245), .Y(n803) );
  OAI21X1 U250 ( .A(n2269), .B(n2305), .C(n1273), .Y(n804) );
  OAI21X1 U252 ( .A(n2268), .B(n2305), .C(n84), .Y(n805) );
  OAI21X1 U254 ( .A(n2267), .B(n2305), .C(n280), .Y(n806) );
  OAI21X1 U256 ( .A(n2266), .B(n2305), .C(n1496), .Y(n807) );
  OAI21X1 U258 ( .A(n2265), .B(n2305), .C(n1532), .Y(n808) );
  OAI21X1 U260 ( .A(n2264), .B(n2305), .C(n1363), .Y(n809) );
  OAI21X1 U262 ( .A(n2263), .B(n2305), .C(n1395), .Y(n810) );
  OAI21X1 U265 ( .A(n2278), .B(n2304), .C(n1462), .Y(n811) );
  OAI21X1 U267 ( .A(n2277), .B(n2304), .C(n1428), .Y(n812) );
  OAI21X1 U269 ( .A(n2276), .B(n2304), .C(n1531), .Y(n813) );
  OAI21X1 U271 ( .A(n2275), .B(n2304), .C(n1495), .Y(n814) );
  OAI21X1 U273 ( .A(n2274), .B(n2304), .C(n1614), .Y(n815) );
  OAI21X1 U275 ( .A(n2273), .B(n2304), .C(n1573), .Y(n816) );
  OAI21X1 U277 ( .A(n2272), .B(n2304), .C(n1698), .Y(n817) );
  OAI21X1 U279 ( .A(n2271), .B(n2304), .C(n1655), .Y(n818) );
  OAI21X1 U281 ( .A(n2270), .B(n2304), .C(n263), .Y(n819) );
  OAI21X1 U283 ( .A(n2269), .B(n2304), .C(n83), .Y(n820) );
  OAI21X1 U285 ( .A(n2268), .B(n2304), .C(n1272), .Y(n821) );
  OAI21X1 U287 ( .A(n2267), .B(n2304), .C(n1244), .Y(n822) );
  OAI21X1 U289 ( .A(n2266), .B(n2304), .C(n1461), .Y(n823) );
  OAI21X1 U291 ( .A(n2265), .B(n2304), .C(n1427), .Y(n824) );
  OAI21X1 U293 ( .A(n2264), .B(n2304), .C(n1332), .Y(n825) );
  OAI21X1 U295 ( .A(n2263), .B(n2304), .C(n1302), .Y(n826) );
  OAI21X1 U298 ( .A(n2278), .B(n2303), .C(n1426), .Y(n827) );
  OAI21X1 U300 ( .A(n2277), .B(n2303), .C(n1460), .Y(n828) );
  OAI21X1 U302 ( .A(n2276), .B(n2303), .C(n1494), .Y(n829) );
  OAI21X1 U304 ( .A(n2275), .B(n2303), .C(n1530), .Y(n830) );
  OAI21X1 U306 ( .A(n2274), .B(n2303), .C(n1572), .Y(n831) );
  OAI21X1 U308 ( .A(n2273), .B(n2303), .C(n1613), .Y(n832) );
  OAI21X1 U310 ( .A(n2272), .B(n2303), .C(n1654), .Y(n833) );
  OAI21X1 U312 ( .A(n2271), .B(n2303), .C(n1697), .Y(n834) );
  OAI21X1 U314 ( .A(n2270), .B(n2303), .C(n76), .Y(n835) );
  OAI21X1 U316 ( .A(n2269), .B(n2303), .C(n245), .Y(n836) );
  OAI21X1 U318 ( .A(n2268), .B(n2303), .C(n1243), .Y(n837) );
  OAI21X1 U320 ( .A(n2267), .B(n2303), .C(n1271), .Y(n838) );
  OAI21X1 U322 ( .A(n2266), .B(n2303), .C(n1425), .Y(n839) );
  OAI21X1 U324 ( .A(n2265), .B(n2303), .C(n1459), .Y(n840) );
  OAI21X1 U326 ( .A(n2264), .B(n2303), .C(n1301), .Y(n841) );
  OAI21X1 U328 ( .A(n2263), .B(n2303), .C(n1331), .Y(n842) );
  NOR3X1 U331 ( .A(wr_ptr[3]), .B(wr_ptr[4]), .C(n658), .Y(n118) );
  OAI21X1 U332 ( .A(n2278), .B(n2302), .C(n1394), .Y(n843) );
  OAI21X1 U334 ( .A(n2277), .B(n2302), .C(n1362), .Y(n844) );
  OAI21X1 U336 ( .A(n2276), .B(n2302), .C(n1330), .Y(n845) );
  OAI21X1 U338 ( .A(n2275), .B(n2302), .C(n1300), .Y(n846) );
  OAI21X1 U340 ( .A(n2274), .B(n2302), .C(n1270), .Y(n847) );
  OAI21X1 U342 ( .A(n2273), .B(n2302), .C(n1242), .Y(n848) );
  OAI21X1 U344 ( .A(n2272), .B(n2302), .C(n227), .Y(n849) );
  OAI21X1 U346 ( .A(n2271), .B(n2302), .C(n75), .Y(n850) );
  OAI21X1 U348 ( .A(n2270), .B(n2302), .C(n1696), .Y(n851) );
  OAI21X1 U350 ( .A(n2269), .B(n2302), .C(n1653), .Y(n852) );
  OAI21X1 U352 ( .A(n2268), .B(n2302), .C(n1612), .Y(n853) );
  OAI21X1 U354 ( .A(n2267), .B(n2302), .C(n1571), .Y(n854) );
  OAI21X1 U356 ( .A(n2266), .B(n2302), .C(n1393), .Y(n855) );
  OAI21X1 U358 ( .A(n2265), .B(n2302), .C(n1361), .Y(n856) );
  OAI21X1 U360 ( .A(n2264), .B(n2302), .C(n1529), .Y(n857) );
  OAI21X1 U362 ( .A(n2263), .B(n2302), .C(n1493), .Y(n858) );
  OAI21X1 U365 ( .A(n2278), .B(n2301), .C(n1360), .Y(n859) );
  OAI21X1 U367 ( .A(n2277), .B(n2301), .C(n1392), .Y(n860) );
  OAI21X1 U369 ( .A(n2276), .B(n2301), .C(n1299), .Y(n861) );
  OAI21X1 U371 ( .A(n2275), .B(n2301), .C(n1329), .Y(n862) );
  OAI21X1 U373 ( .A(n2274), .B(n2301), .C(n1241), .Y(n863) );
  OAI21X1 U375 ( .A(n2273), .B(n2301), .C(n1269), .Y(n864) );
  OAI21X1 U377 ( .A(n2272), .B(n2301), .C(n74), .Y(n865) );
  OAI21X1 U379 ( .A(n2271), .B(n2301), .C(n209), .Y(n866) );
  OAI21X1 U381 ( .A(n2270), .B(n2301), .C(n1652), .Y(n867) );
  OAI21X1 U383 ( .A(n2269), .B(n2301), .C(n1695), .Y(n868) );
  OAI21X1 U385 ( .A(n2268), .B(n2301), .C(n1570), .Y(n869) );
  OAI21X1 U387 ( .A(n2267), .B(n2301), .C(n1611), .Y(n870) );
  OAI21X1 U389 ( .A(n2266), .B(n2301), .C(n1359), .Y(n871) );
  OAI21X1 U391 ( .A(n2265), .B(n2301), .C(n1391), .Y(n872) );
  OAI21X1 U393 ( .A(n2264), .B(n2301), .C(n1492), .Y(n873) );
  OAI21X1 U395 ( .A(n2263), .B(n2301), .C(n1528), .Y(n874) );
  OAI21X1 U398 ( .A(n2278), .B(n2300), .C(n1328), .Y(n875) );
  OAI21X1 U400 ( .A(n2277), .B(n2300), .C(n1298), .Y(n876) );
  OAI21X1 U402 ( .A(n2276), .B(n2300), .C(n1390), .Y(n877) );
  OAI21X1 U404 ( .A(n2275), .B(n2300), .C(n1358), .Y(n878) );
  OAI21X1 U406 ( .A(n2274), .B(n2300), .C(n191), .Y(n879) );
  OAI21X1 U408 ( .A(n2273), .B(n2300), .C(n73), .Y(n880) );
  OAI21X1 U410 ( .A(n2272), .B(n2300), .C(n1268), .Y(n881) );
  OAI21X1 U412 ( .A(n2271), .B(n2300), .C(n1240), .Y(n882) );
  OAI21X1 U414 ( .A(n2270), .B(n2300), .C(n1610), .Y(n883) );
  OAI21X1 U416 ( .A(n2269), .B(n2300), .C(n1569), .Y(n884) );
  OAI21X1 U418 ( .A(n2268), .B(n2300), .C(n1694), .Y(n885) );
  OAI21X1 U420 ( .A(n2267), .B(n2300), .C(n1651), .Y(n886) );
  OAI21X1 U422 ( .A(n2266), .B(n2300), .C(n1327), .Y(n887) );
  OAI21X1 U424 ( .A(n2265), .B(n2300), .C(n1297), .Y(n888) );
  OAI21X1 U426 ( .A(n2264), .B(n2300), .C(n1458), .Y(n889) );
  OAI21X1 U428 ( .A(n2263), .B(n2300), .C(n1424), .Y(n890) );
  OAI21X1 U431 ( .A(n2278), .B(n2299), .C(n1296), .Y(n891) );
  OAI21X1 U433 ( .A(n2277), .B(n2299), .C(n1326), .Y(n892) );
  OAI21X1 U435 ( .A(n2276), .B(n2299), .C(n1357), .Y(n893) );
  OAI21X1 U437 ( .A(n2275), .B(n2299), .C(n1389), .Y(n894) );
  OAI21X1 U439 ( .A(n2274), .B(n2299), .C(n72), .Y(n895) );
  OAI21X1 U441 ( .A(n2273), .B(n2299), .C(n173), .Y(n896) );
  OAI21X1 U443 ( .A(n2272), .B(n2299), .C(n666), .Y(n897) );
  OAI21X1 U445 ( .A(n2271), .B(n2299), .C(n1267), .Y(n898) );
  OAI21X1 U447 ( .A(n2270), .B(n2299), .C(n1568), .Y(n899) );
  OAI21X1 U449 ( .A(n2269), .B(n2299), .C(n1609), .Y(n900) );
  OAI21X1 U451 ( .A(n2268), .B(n2299), .C(n1650), .Y(n901) );
  OAI21X1 U453 ( .A(n2267), .B(n2299), .C(n1693), .Y(n902) );
  OAI21X1 U455 ( .A(n2266), .B(n2299), .C(n1295), .Y(n903) );
  OAI21X1 U457 ( .A(n2265), .B(n2299), .C(n1325), .Y(n904) );
  OAI21X1 U459 ( .A(n2264), .B(n2299), .C(n1423), .Y(n905) );
  OAI21X1 U461 ( .A(n2263), .B(n2299), .C(n1457), .Y(n906) );
  OAI21X1 U464 ( .A(n2278), .B(n2298), .C(n1266), .Y(n907) );
  OAI21X1 U466 ( .A(n2277), .B(n2298), .C(n639), .Y(n908) );
  OAI21X1 U468 ( .A(n2276), .B(n2298), .C(n155), .Y(n909) );
  OAI21X1 U470 ( .A(n2275), .B(n2298), .C(n71), .Y(n910) );
  OAI21X1 U472 ( .A(n2274), .B(n2298), .C(n1388), .Y(n911) );
  OAI21X1 U474 ( .A(n2273), .B(n2298), .C(n1356), .Y(n912) );
  OAI21X1 U476 ( .A(n2272), .B(n2298), .C(n1324), .Y(n913) );
  OAI21X1 U478 ( .A(n2271), .B(n2298), .C(n1294), .Y(n914) );
  OAI21X1 U480 ( .A(n2270), .B(n2298), .C(n1527), .Y(n915) );
  OAI21X1 U482 ( .A(n2269), .B(n2298), .C(n1491), .Y(n916) );
  OAI21X1 U484 ( .A(n2268), .B(n2298), .C(n1456), .Y(n917) );
  OAI21X1 U486 ( .A(n2267), .B(n2298), .C(n1422), .Y(n918) );
  OAI21X1 U488 ( .A(n2266), .B(n2298), .C(n1265), .Y(n919) );
  OAI21X1 U490 ( .A(n2265), .B(n2298), .C(n622), .Y(n920) );
  OAI21X1 U492 ( .A(n2264), .B(n2298), .C(n1692), .Y(n921) );
  OAI21X1 U494 ( .A(n2263), .B(n2298), .C(n1649), .Y(n922) );
  OAI21X1 U497 ( .A(n2278), .B(n2297), .C(n1691), .Y(n923) );
  OAI21X1 U499 ( .A(n2277), .B(n2297), .C(n1648), .Y(n924) );
  OAI21X1 U501 ( .A(n2276), .B(n2297), .C(n1608), .Y(n925) );
  OAI21X1 U503 ( .A(n2275), .B(n2297), .C(n1567), .Y(n926) );
  OAI21X1 U505 ( .A(n2274), .B(n2297), .C(n1526), .Y(n927) );
  OAI21X1 U507 ( .A(n2273), .B(n2297), .C(n1490), .Y(n928) );
  OAI21X1 U509 ( .A(n2272), .B(n2297), .C(n1455), .Y(n929) );
  OAI21X1 U511 ( .A(n2271), .B(n2297), .C(n1421), .Y(n930) );
  OAI21X1 U513 ( .A(n2270), .B(n2297), .C(n1387), .Y(n931) );
  OAI21X1 U515 ( .A(n2269), .B(n2297), .C(n1355), .Y(n932) );
  OAI21X1 U517 ( .A(n2268), .B(n2297), .C(n1323), .Y(n933) );
  OAI21X1 U519 ( .A(n2267), .B(n2297), .C(n1293), .Y(n934) );
  OAI21X1 U521 ( .A(n2266), .B(n2297), .C(n1690), .Y(n935) );
  OAI21X1 U523 ( .A(n2265), .B(n2297), .C(n1647), .Y(n936) );
  OAI21X1 U525 ( .A(n2264), .B(n2297), .C(n1264), .Y(n937) );
  OAI21X1 U527 ( .A(n2263), .B(n2297), .C(n605), .Y(n938) );
  OAI21X1 U530 ( .A(n2278), .B(n2296), .C(n1646), .Y(n939) );
  OAI21X1 U532 ( .A(n2277), .B(n2296), .C(n1689), .Y(n940) );
  OAI21X1 U534 ( .A(n2276), .B(n2296), .C(n1566), .Y(n941) );
  OAI21X1 U536 ( .A(n2275), .B(n2296), .C(n1607), .Y(n942) );
  OAI21X1 U538 ( .A(n2274), .B(n2296), .C(n1489), .Y(n943) );
  OAI21X1 U540 ( .A(n2273), .B(n2296), .C(n1525), .Y(n944) );
  OAI21X1 U542 ( .A(n2272), .B(n2296), .C(n1420), .Y(n945) );
  OAI21X1 U544 ( .A(n2271), .B(n2296), .C(n1454), .Y(n946) );
  OAI21X1 U546 ( .A(n2270), .B(n2296), .C(n1354), .Y(n947) );
  OAI21X1 U548 ( .A(n2269), .B(n2296), .C(n1386), .Y(n948) );
  OAI21X1 U550 ( .A(n2268), .B(n2296), .C(n1292), .Y(n949) );
  OAI21X1 U552 ( .A(n2267), .B(n2296), .C(n1322), .Y(n950) );
  OAI21X1 U554 ( .A(n2266), .B(n2296), .C(n1645), .Y(n951) );
  OAI21X1 U556 ( .A(n2265), .B(n2296), .C(n1688), .Y(n952) );
  OAI21X1 U558 ( .A(n2264), .B(n2296), .C(n588), .Y(n953) );
  OAI21X1 U560 ( .A(n2263), .B(n2296), .C(n1263), .Y(n954) );
  OAI21X1 U563 ( .A(n2278), .B(n2295), .C(n1606), .Y(n955) );
  OAI21X1 U565 ( .A(n2277), .B(n2295), .C(n1565), .Y(n956) );
  OAI21X1 U567 ( .A(n2276), .B(n2295), .C(n1687), .Y(n957) );
  OAI21X1 U569 ( .A(n2275), .B(n2295), .C(n1644), .Y(n958) );
  OAI21X1 U571 ( .A(n2274), .B(n2295), .C(n1453), .Y(n959) );
  OAI21X1 U573 ( .A(n2273), .B(n2295), .C(n1419), .Y(n960) );
  OAI21X1 U575 ( .A(n2272), .B(n2295), .C(n1524), .Y(n961) );
  OAI21X1 U577 ( .A(n2271), .B(n2295), .C(n1488), .Y(n962) );
  OAI21X1 U579 ( .A(n2270), .B(n2295), .C(n1321), .Y(n963) );
  OAI21X1 U581 ( .A(n2269), .B(n2295), .C(n1291), .Y(n964) );
  OAI21X1 U583 ( .A(n2268), .B(n2295), .C(n1385), .Y(n965) );
  OAI21X1 U585 ( .A(n2267), .B(n2295), .C(n1353), .Y(n966) );
  OAI21X1 U587 ( .A(n2266), .B(n2295), .C(n1605), .Y(n967) );
  OAI21X1 U589 ( .A(n2265), .B(n2295), .C(n1564), .Y(n968) );
  OAI21X1 U591 ( .A(n2264), .B(n2295), .C(n137), .Y(n969) );
  OAI21X1 U593 ( .A(n2263), .B(n2295), .C(n65), .Y(n970) );
  NOR3X1 U596 ( .A(n658), .B(wr_ptr[4]), .C(n2347), .Y(n262) );
  OAI21X1 U597 ( .A(n2278), .B(n2294), .C(n1563), .Y(n971) );
  OAI21X1 U599 ( .A(n2277), .B(n2294), .C(n1604), .Y(n972) );
  OAI21X1 U601 ( .A(n2276), .B(n2294), .C(n1643), .Y(n973) );
  OAI21X1 U603 ( .A(n2275), .B(n2294), .C(n1686), .Y(n974) );
  OAI21X1 U605 ( .A(n2274), .B(n2294), .C(n1418), .Y(n975) );
  OAI21X1 U607 ( .A(n2273), .B(n2294), .C(n1452), .Y(n976) );
  OAI21X1 U609 ( .A(n2272), .B(n2294), .C(n1487), .Y(n977) );
  OAI21X1 U611 ( .A(n2271), .B(n2294), .C(n1523), .Y(n978) );
  OAI21X1 U613 ( .A(n2270), .B(n2294), .C(n1290), .Y(n979) );
  OAI21X1 U615 ( .A(n2269), .B(n2294), .C(n1320), .Y(n980) );
  OAI21X1 U617 ( .A(n2268), .B(n2294), .C(n1352), .Y(n981) );
  OAI21X1 U619 ( .A(n2267), .B(n2294), .C(n1384), .Y(n982) );
  OAI21X1 U621 ( .A(n2266), .B(n2294), .C(n1562), .Y(n983) );
  OAI21X1 U623 ( .A(n2265), .B(n2294), .C(n1603), .Y(n984) );
  OAI21X1 U625 ( .A(n2264), .B(n2294), .C(n64), .Y(n985) );
  OAI21X1 U627 ( .A(n2263), .B(n2294), .C(n119), .Y(n986) );
  OAI21X1 U630 ( .A(n2278), .B(n2293), .C(n1522), .Y(n987) );
  OAI21X1 U632 ( .A(n2277), .B(n2293), .C(n1486), .Y(n988) );
  OAI21X1 U634 ( .A(n2276), .B(n2293), .C(n1451), .Y(n989) );
  OAI21X1 U636 ( .A(n2275), .B(n2293), .C(n1417), .Y(n990) );
  OAI21X1 U638 ( .A(n2274), .B(n2293), .C(n1685), .Y(n991) );
  OAI21X1 U640 ( .A(n2273), .B(n2293), .C(n1642), .Y(n992) );
  OAI21X1 U642 ( .A(n2272), .B(n2293), .C(n1602), .Y(n993) );
  OAI21X1 U644 ( .A(n2271), .B(n2293), .C(n1561), .Y(n994) );
  OAI21X1 U646 ( .A(n2270), .B(n2293), .C(n1262), .Y(n995) );
  OAI21X1 U648 ( .A(n2269), .B(n2293), .C(n571), .Y(n996) );
  OAI21X1 U650 ( .A(n2268), .B(n2293), .C(n100), .Y(n997) );
  OAI21X1 U652 ( .A(n2267), .B(n2293), .C(n63), .Y(n998) );
  OAI21X1 U654 ( .A(n2266), .B(n2293), .C(n1521), .Y(n999) );
  OAI21X1 U656 ( .A(n2265), .B(n2293), .C(n1485), .Y(n1000) );
  OAI21X1 U658 ( .A(n2264), .B(n2293), .C(n1383), .Y(n1001) );
  OAI21X1 U660 ( .A(n2263), .B(n2293), .C(n1351), .Y(n1002) );
  OAI21X1 U663 ( .A(n2278), .B(n2292), .C(n1484), .Y(n1003) );
  OAI21X1 U665 ( .A(n2277), .B(n2292), .C(n1520), .Y(n1004) );
  OAI21X1 U667 ( .A(n2276), .B(n2292), .C(n1416), .Y(n1005) );
  OAI21X1 U669 ( .A(n2275), .B(n2292), .C(n1450), .Y(n1006) );
  OAI21X1 U671 ( .A(n2274), .B(n2292), .C(n1641), .Y(n1007) );
  OAI21X1 U673 ( .A(n2273), .B(n2292), .C(n1684), .Y(n1008) );
  OAI21X1 U675 ( .A(n2272), .B(n2292), .C(n1560), .Y(n1009) );
  OAI21X1 U677 ( .A(n2271), .B(n2292), .C(n1601), .Y(n1010) );
  OAI21X1 U679 ( .A(n2270), .B(n2292), .C(n554), .Y(n1011) );
  OAI21X1 U681 ( .A(n2269), .B(n2292), .C(n1261), .Y(n1012) );
  OAI21X1 U683 ( .A(n2268), .B(n2292), .C(n62), .Y(n1013) );
  OAI21X1 U685 ( .A(n2267), .B(n2292), .C(n99), .Y(n1014) );
  OAI21X1 U687 ( .A(n2266), .B(n2292), .C(n1483), .Y(n1015) );
  OAI21X1 U689 ( .A(n2265), .B(n2292), .C(n1519), .Y(n1016) );
  OAI21X1 U691 ( .A(n2264), .B(n2292), .C(n1350), .Y(n1017) );
  OAI21X1 U693 ( .A(n2263), .B(n2292), .C(n1382), .Y(n1018) );
  OAI21X1 U696 ( .A(n2278), .B(n2291), .C(n1449), .Y(n1019) );
  OAI21X1 U698 ( .A(n2277), .B(n2291), .C(n1415), .Y(n1020) );
  OAI21X1 U700 ( .A(n2276), .B(n2291), .C(n1518), .Y(n1021) );
  OAI21X1 U702 ( .A(n2275), .B(n2291), .C(n1482), .Y(n1022) );
  OAI21X1 U704 ( .A(n2274), .B(n2291), .C(n1600), .Y(n1023) );
  OAI21X1 U706 ( .A(n2273), .B(n2291), .C(n1559), .Y(n1024) );
  OAI21X1 U708 ( .A(n2272), .B(n2291), .C(n1683), .Y(n1025) );
  OAI21X1 U710 ( .A(n2271), .B(n2291), .C(n1640), .Y(n1026) );
  OAI21X1 U712 ( .A(n2270), .B(n2291), .C(n98), .Y(n1027) );
  OAI21X1 U714 ( .A(n2269), .B(n2291), .C(n61), .Y(n1028) );
  OAI21X1 U716 ( .A(n2268), .B(n2291), .C(n1260), .Y(n1029) );
  OAI21X1 U718 ( .A(n2267), .B(n2291), .C(n537), .Y(n1030) );
  OAI21X1 U720 ( .A(n2266), .B(n2291), .C(n1448), .Y(n1031) );
  OAI21X1 U722 ( .A(n2265), .B(n2291), .C(n1414), .Y(n1032) );
  OAI21X1 U724 ( .A(n2264), .B(n2291), .C(n1319), .Y(n1033) );
  OAI21X1 U726 ( .A(n2263), .B(n2291), .C(n1289), .Y(n1034) );
  OAI21X1 U729 ( .A(n2278), .B(n2290), .C(n1413), .Y(n1035) );
  OAI21X1 U731 ( .A(n2277), .B(n2290), .C(n1447), .Y(n1036) );
  OAI21X1 U733 ( .A(n2276), .B(n2290), .C(n1481), .Y(n1037) );
  OAI21X1 U735 ( .A(n2275), .B(n2290), .C(n1517), .Y(n1038) );
  OAI21X1 U737 ( .A(n2274), .B(n2290), .C(n1558), .Y(n1039) );
  OAI21X1 U739 ( .A(n2273), .B(n2290), .C(n1599), .Y(n1040) );
  OAI21X1 U741 ( .A(n2272), .B(n2290), .C(n1639), .Y(n1041) );
  OAI21X1 U743 ( .A(n2271), .B(n2290), .C(n1682), .Y(n1042) );
  OAI21X1 U745 ( .A(n2270), .B(n2290), .C(n60), .Y(n1043) );
  OAI21X1 U747 ( .A(n2269), .B(n2290), .C(n97), .Y(n1044) );
  OAI21X1 U749 ( .A(n2268), .B(n2290), .C(n519), .Y(n1045) );
  OAI21X1 U751 ( .A(n2267), .B(n2290), .C(n1259), .Y(n1046) );
  OAI21X1 U753 ( .A(n2266), .B(n2290), .C(n1412), .Y(n1047) );
  OAI21X1 U755 ( .A(n2265), .B(n2290), .C(n1446), .Y(n1048) );
  OAI21X1 U757 ( .A(n2264), .B(n2290), .C(n1288), .Y(n1049) );
  OAI21X1 U759 ( .A(n2263), .B(n2290), .C(n1318), .Y(n1050) );
  OAI21X1 U762 ( .A(n2278), .B(n2289), .C(n1381), .Y(n1051) );
  OAI21X1 U764 ( .A(n2277), .B(n2289), .C(n1349), .Y(n1052) );
  OAI21X1 U766 ( .A(n2276), .B(n2289), .C(n1317), .Y(n1053) );
  OAI21X1 U768 ( .A(n2275), .B(n2289), .C(n1287), .Y(n1054) );
  OAI21X1 U770 ( .A(n2274), .B(n2289), .C(n1258), .Y(n1055) );
  OAI21X1 U772 ( .A(n2273), .B(n2289), .C(n502), .Y(n1056) );
  OAI21X1 U774 ( .A(n2272), .B(n2289), .C(n96), .Y(n1057) );
  OAI21X1 U776 ( .A(n2271), .B(n2289), .C(n59), .Y(n1058) );
  OAI21X1 U778 ( .A(n2270), .B(n2289), .C(n1681), .Y(n1059) );
  OAI21X1 U780 ( .A(n2269), .B(n2289), .C(n1638), .Y(n1060) );
  OAI21X1 U782 ( .A(n2268), .B(n2289), .C(n1598), .Y(n1061) );
  OAI21X1 U784 ( .A(n2267), .B(n2289), .C(n1557), .Y(n1062) );
  OAI21X1 U786 ( .A(n2266), .B(n2289), .C(n1380), .Y(n1063) );
  OAI21X1 U788 ( .A(n2265), .B(n2289), .C(n1348), .Y(n1064) );
  OAI21X1 U790 ( .A(n2264), .B(n2289), .C(n1516), .Y(n1065) );
  OAI21X1 U792 ( .A(n2263), .B(n2289), .C(n1480), .Y(n1066) );
  OAI21X1 U795 ( .A(n2278), .B(n2288), .C(n1347), .Y(n1067) );
  OAI21X1 U797 ( .A(n2277), .B(n2288), .C(n1379), .Y(n1068) );
  OAI21X1 U799 ( .A(n2276), .B(n2288), .C(n1286), .Y(n1069) );
  OAI21X1 U801 ( .A(n2275), .B(n2288), .C(n1316), .Y(n1070) );
  OAI21X1 U803 ( .A(n2274), .B(n2288), .C(n485), .Y(n1071) );
  OAI21X1 U805 ( .A(n2273), .B(n2288), .C(n1257), .Y(n1072) );
  OAI21X1 U807 ( .A(n2272), .B(n2288), .C(n54), .Y(n1073) );
  OAI21X1 U809 ( .A(n2271), .B(n2288), .C(n95), .Y(n1074) );
  OAI21X1 U811 ( .A(n2270), .B(n2288), .C(n1637), .Y(n1075) );
  OAI21X1 U813 ( .A(n2269), .B(n2288), .C(n1680), .Y(n1076) );
  OAI21X1 U815 ( .A(n2268), .B(n2288), .C(n1556), .Y(n1077) );
  OAI21X1 U817 ( .A(n2267), .B(n2288), .C(n1597), .Y(n1078) );
  OAI21X1 U819 ( .A(n2266), .B(n2288), .C(n1346), .Y(n1079) );
  OAI21X1 U821 ( .A(n2265), .B(n2288), .C(n1378), .Y(n1080) );
  OAI21X1 U823 ( .A(n2264), .B(n2288), .C(n1479), .Y(n1081) );
  OAI21X1 U825 ( .A(n2263), .B(n2288), .C(n1515), .Y(n1082) );
  OAI21X1 U828 ( .A(n2278), .B(n2287), .C(n1315), .Y(n1083) );
  OAI21X1 U830 ( .A(n2277), .B(n2287), .C(n1285), .Y(n1084) );
  OAI21X1 U832 ( .A(n2276), .B(n2287), .C(n1377), .Y(n1085) );
  OAI21X1 U834 ( .A(n2275), .B(n2287), .C(n1345), .Y(n1086) );
  OAI21X1 U836 ( .A(n2274), .B(n2287), .C(n94), .Y(n1087) );
  OAI21X1 U838 ( .A(n2273), .B(n2287), .C(n49), .Y(n1088) );
  OAI21X1 U840 ( .A(n2272), .B(n2287), .C(n1256), .Y(n1089) );
  OAI21X1 U842 ( .A(n2271), .B(n2287), .C(n468), .Y(n1090) );
  OAI21X1 U844 ( .A(n2270), .B(n2287), .C(n1596), .Y(n1091) );
  OAI21X1 U846 ( .A(n2269), .B(n2287), .C(n1555), .Y(n1092) );
  OAI21X1 U848 ( .A(n2268), .B(n2287), .C(n1679), .Y(n1093) );
  OAI21X1 U850 ( .A(n2267), .B(n2287), .C(n1636), .Y(n1094) );
  OAI21X1 U852 ( .A(n2266), .B(n2287), .C(n1314), .Y(n1095) );
  OAI21X1 U854 ( .A(n2265), .B(n2287), .C(n1284), .Y(n1096) );
  OAI21X1 U856 ( .A(n2264), .B(n2287), .C(n1445), .Y(n1097) );
  OAI21X1 U858 ( .A(n2263), .B(n2287), .C(n1411), .Y(n1098) );
  NOR3X1 U861 ( .A(n658), .B(wr_ptr[3]), .C(n2348), .Y(n399) );
  OAI21X1 U862 ( .A(n2278), .B(n2286), .C(n1283), .Y(n1099) );
  OAI21X1 U864 ( .A(n2277), .B(n2286), .C(n1313), .Y(n1100) );
  OAI21X1 U866 ( .A(n2276), .B(n2286), .C(n1344), .Y(n1101) );
  OAI21X1 U868 ( .A(n2275), .B(n2286), .C(n1376), .Y(n1102) );
  OAI21X1 U870 ( .A(n2274), .B(n2286), .C(n48), .Y(n1103) );
  OAI21X1 U872 ( .A(n2273), .B(n2286), .C(n93), .Y(n1104) );
  OAI21X1 U874 ( .A(n2272), .B(n2286), .C(n451), .Y(n1105) );
  OAI21X1 U876 ( .A(n2271), .B(n2286), .C(n1255), .Y(n1106) );
  OAI21X1 U878 ( .A(n2270), .B(n2286), .C(n1554), .Y(n1107) );
  OAI21X1 U880 ( .A(n2269), .B(n2286), .C(n1595), .Y(n1108) );
  OAI21X1 U882 ( .A(n2268), .B(n2286), .C(n1635), .Y(n1109) );
  OAI21X1 U884 ( .A(n2267), .B(n2286), .C(n1678), .Y(n1110) );
  OAI21X1 U886 ( .A(n2266), .B(n2286), .C(n1282), .Y(n1111) );
  OAI21X1 U888 ( .A(n2265), .B(n2286), .C(n1312), .Y(n1112) );
  OAI21X1 U890 ( .A(n2264), .B(n2286), .C(n1410), .Y(n1113) );
  OAI21X1 U892 ( .A(n2263), .B(n2286), .C(n1444), .Y(n1114) );
  NOR3X1 U895 ( .A(wr_ptr[1]), .B(wr_ptr[2]), .C(wr_ptr[0]), .Y(n117) );
  OAI21X1 U896 ( .A(n2278), .B(n2285), .C(n1254), .Y(n1115) );
  OAI21X1 U898 ( .A(n2277), .B(n2285), .C(n434), .Y(n1116) );
  OAI21X1 U900 ( .A(n2276), .B(n2285), .C(n92), .Y(n1117) );
  OAI21X1 U902 ( .A(n2275), .B(n2285), .C(n47), .Y(n1118) );
  OAI21X1 U904 ( .A(n2274), .B(n2285), .C(n1375), .Y(n1119) );
  OAI21X1 U906 ( .A(n2273), .B(n2285), .C(n1343), .Y(n1120) );
  OAI21X1 U908 ( .A(n2272), .B(n2285), .C(n1311), .Y(n1121) );
  OAI21X1 U910 ( .A(n2271), .B(n2285), .C(n1281), .Y(n1122) );
  OAI21X1 U912 ( .A(n2270), .B(n2285), .C(n1514), .Y(n1123) );
  OAI21X1 U914 ( .A(n2269), .B(n2285), .C(n1478), .Y(n1124) );
  OAI21X1 U916 ( .A(n2268), .B(n2285), .C(n1443), .Y(n1125) );
  OAI21X1 U918 ( .A(n2267), .B(n2285), .C(n1409), .Y(n1126) );
  OAI21X1 U920 ( .A(n2266), .B(n2285), .C(n1253), .Y(n1127) );
  OAI21X1 U922 ( .A(n2265), .B(n2285), .C(n417), .Y(n1128) );
  OAI21X1 U924 ( .A(n2264), .B(n2285), .C(n1677), .Y(n1129) );
  OAI21X1 U926 ( .A(n2263), .B(n2285), .C(n1634), .Y(n1130) );
  NOR3X1 U929 ( .A(wr_ptr[1]), .B(wr_ptr[2]), .C(n2344), .Y(n136) );
  OAI21X1 U930 ( .A(n2278), .B(n2284), .C(n1676), .Y(n1131) );
  OAI21X1 U932 ( .A(n2277), .B(n2284), .C(n1633), .Y(n1132) );
  OAI21X1 U934 ( .A(n2276), .B(n2284), .C(n1594), .Y(n1133) );
  OAI21X1 U936 ( .A(n2275), .B(n2284), .C(n1553), .Y(n1134) );
  OAI21X1 U938 ( .A(n2274), .B(n2284), .C(n1513), .Y(n1135) );
  OAI21X1 U940 ( .A(n2273), .B(n2284), .C(n1477), .Y(n1136) );
  OAI21X1 U942 ( .A(n2272), .B(n2284), .C(n1442), .Y(n1137) );
  OAI21X1 U944 ( .A(n2271), .B(n2284), .C(n1408), .Y(n1138) );
  OAI21X1 U946 ( .A(n2270), .B(n2284), .C(n1374), .Y(n1139) );
  OAI21X1 U948 ( .A(n2269), .B(n2284), .C(n1342), .Y(n1140) );
  OAI21X1 U950 ( .A(n2268), .B(n2284), .C(n1310), .Y(n1141) );
  OAI21X1 U952 ( .A(n2267), .B(n2284), .C(n1280), .Y(n1142) );
  OAI21X1 U954 ( .A(n2266), .B(n2284), .C(n1675), .Y(n1143) );
  OAI21X1 U956 ( .A(n2265), .B(n2284), .C(n1632), .Y(n1144) );
  OAI21X1 U958 ( .A(n2264), .B(n2284), .C(n1252), .Y(n1145) );
  OAI21X1 U960 ( .A(n2263), .B(n2284), .C(n400), .Y(n1146) );
  NOR3X1 U963 ( .A(wr_ptr[0]), .B(wr_ptr[2]), .C(n2345), .Y(n154) );
  OAI21X1 U964 ( .A(n2278), .B(n2283), .C(n1631), .Y(n1147) );
  OAI21X1 U966 ( .A(n2277), .B(n2283), .C(n1674), .Y(n1148) );
  OAI21X1 U968 ( .A(n2276), .B(n2283), .C(n1552), .Y(n1149) );
  OAI21X1 U970 ( .A(n2275), .B(n2283), .C(n1593), .Y(n1150) );
  OAI21X1 U972 ( .A(n2274), .B(n2283), .C(n1476), .Y(n1151) );
  OAI21X1 U974 ( .A(n2273), .B(n2283), .C(n1512), .Y(n1152) );
  OAI21X1 U976 ( .A(n2272), .B(n2283), .C(n1407), .Y(n1153) );
  OAI21X1 U978 ( .A(n2271), .B(n2283), .C(n1441), .Y(n1154) );
  OAI21X1 U980 ( .A(n2270), .B(n2283), .C(n1341), .Y(n1155) );
  OAI21X1 U982 ( .A(n2269), .B(n2283), .C(n1373), .Y(n1156) );
  OAI21X1 U984 ( .A(n2268), .B(n2283), .C(n1279), .Y(n1157) );
  OAI21X1 U986 ( .A(n2267), .B(n2283), .C(n1309), .Y(n1158) );
  OAI21X1 U988 ( .A(n2266), .B(n2283), .C(n1630), .Y(n1159) );
  OAI21X1 U990 ( .A(n2265), .B(n2283), .C(n1673), .Y(n1160) );
  OAI21X1 U992 ( .A(n2264), .B(n2283), .C(n382), .Y(n1161) );
  OAI21X1 U994 ( .A(n2263), .B(n2283), .C(n1251), .Y(n1162) );
  NOR3X1 U997 ( .A(n2344), .B(wr_ptr[2]), .C(n2345), .Y(n172) );
  OAI21X1 U998 ( .A(n2278), .B(n2282), .C(n1592), .Y(n1163) );
  OAI21X1 U1000 ( .A(n2277), .B(n2282), .C(n1551), .Y(n1164) );
  OAI21X1 U1002 ( .A(n2276), .B(n2282), .C(n1672), .Y(n1165) );
  OAI21X1 U1004 ( .A(n2275), .B(n2282), .C(n1629), .Y(n1166) );
  OAI21X1 U1006 ( .A(n2274), .B(n2282), .C(n1440), .Y(n1167) );
  OAI21X1 U1008 ( .A(n2273), .B(n2282), .C(n1406), .Y(n1168) );
  OAI21X1 U1010 ( .A(n2272), .B(n2282), .C(n1511), .Y(n1169) );
  OAI21X1 U1012 ( .A(n2271), .B(n2282), .C(n1475), .Y(n1170) );
  OAI21X1 U1014 ( .A(n2270), .B(n2282), .C(n1308), .Y(n1171) );
  OAI21X1 U1016 ( .A(n2269), .B(n2282), .C(n1278), .Y(n1172) );
  OAI21X1 U1018 ( .A(n2268), .B(n2282), .C(n1372), .Y(n1173) );
  OAI21X1 U1020 ( .A(n2267), .B(n2282), .C(n1340), .Y(n1174) );
  OAI21X1 U1022 ( .A(n2266), .B(n2282), .C(n1591), .Y(n1175) );
  OAI21X1 U1024 ( .A(n2265), .B(n2282), .C(n1550), .Y(n1176) );
  OAI21X1 U1026 ( .A(n2264), .B(n2282), .C(n91), .Y(n1177) );
  OAI21X1 U1028 ( .A(n2263), .B(n2282), .C(n46), .Y(n1178) );
  NOR3X1 U1031 ( .A(wr_ptr[0]), .B(wr_ptr[1]), .C(n2346), .Y(n190) );
  OAI21X1 U1032 ( .A(n2278), .B(n2281), .C(n1549), .Y(n1179) );
  OAI21X1 U1034 ( .A(n2277), .B(n2281), .C(n1590), .Y(n1180) );
  OAI21X1 U1036 ( .A(n2276), .B(n2281), .C(n1628), .Y(n1181) );
  OAI21X1 U1038 ( .A(n2275), .B(n2281), .C(n1671), .Y(n1182) );
  OAI21X1 U1040 ( .A(n2274), .B(n2281), .C(n1405), .Y(n1183) );
  OAI21X1 U1042 ( .A(n2273), .B(n2281), .C(n1439), .Y(n1184) );
  OAI21X1 U1044 ( .A(n2272), .B(n2281), .C(n1474), .Y(n1185) );
  OAI21X1 U1046 ( .A(n2271), .B(n2281), .C(n1510), .Y(n1186) );
  OAI21X1 U1048 ( .A(n2270), .B(n2281), .C(n1277), .Y(n1187) );
  OAI21X1 U1050 ( .A(n2269), .B(n2281), .C(n1307), .Y(n1188) );
  OAI21X1 U1052 ( .A(n2268), .B(n2281), .C(n1339), .Y(n1189) );
  OAI21X1 U1054 ( .A(n2267), .B(n2281), .C(n1371), .Y(n1190) );
  OAI21X1 U1056 ( .A(n2266), .B(n2281), .C(n1548), .Y(n1191) );
  OAI21X1 U1058 ( .A(n2265), .B(n2281), .C(n1589), .Y(n1192) );
  OAI21X1 U1060 ( .A(n2264), .B(n2281), .C(n45), .Y(n1193) );
  OAI21X1 U1062 ( .A(n2263), .B(n2281), .C(n90), .Y(n1194) );
  NOR3X1 U1065 ( .A(n2344), .B(wr_ptr[1]), .C(n2346), .Y(n208) );
  OAI21X1 U1066 ( .A(n2278), .B(n2280), .C(n1509), .Y(n1195) );
  OAI21X1 U1068 ( .A(n2277), .B(n2280), .C(n1473), .Y(n1196) );
  OAI21X1 U1070 ( .A(n2276), .B(n2280), .C(n1438), .Y(n1197) );
  OAI21X1 U1072 ( .A(n2275), .B(n2280), .C(n1404), .Y(n1198) );
  OAI21X1 U1074 ( .A(n2274), .B(n2280), .C(n1670), .Y(n1199) );
  OAI21X1 U1076 ( .A(n2273), .B(n2280), .C(n1627), .Y(n1200) );
  OAI21X1 U1078 ( .A(n2272), .B(n2280), .C(n1588), .Y(n1201) );
  OAI21X1 U1080 ( .A(n2271), .B(n2280), .C(n1547), .Y(n1202) );
  OAI21X1 U1082 ( .A(n2270), .B(n2280), .C(n1250), .Y(n1203) );
  OAI21X1 U1084 ( .A(n2269), .B(n2280), .C(n365), .Y(n1204) );
  OAI21X1 U1086 ( .A(n2268), .B(n2280), .C(n89), .Y(n1205) );
  OAI21X1 U1088 ( .A(n2267), .B(n2280), .C(n44), .Y(n1206) );
  OAI21X1 U1090 ( .A(n2266), .B(n2280), .C(n1508), .Y(n1207) );
  OAI21X1 U1092 ( .A(n2265), .B(n2280), .C(n1472), .Y(n1208) );
  OAI21X1 U1094 ( .A(n2264), .B(n2280), .C(n1370), .Y(n1209) );
  OAI21X1 U1096 ( .A(n2263), .B(n2280), .C(n1338), .Y(n1210) );
  NOR3X1 U1099 ( .A(n2345), .B(wr_ptr[0]), .C(n2346), .Y(n226) );
  OAI21X1 U1100 ( .A(n2278), .B(n2279), .C(n1471), .Y(n1211) );
  OAI21X1 U1102 ( .A(n2277), .B(n2279), .C(n1507), .Y(n1212) );
  OAI21X1 U1104 ( .A(n2276), .B(n2279), .C(n1403), .Y(n1213) );
  OAI21X1 U1106 ( .A(n2275), .B(n2279), .C(n1437), .Y(n1214) );
  OAI21X1 U1108 ( .A(n2274), .B(n2279), .C(n1626), .Y(n1215) );
  OAI21X1 U1110 ( .A(n2273), .B(n2279), .C(n1669), .Y(n1216) );
  OAI21X1 U1112 ( .A(n2272), .B(n2279), .C(n1546), .Y(n1217) );
  OAI21X1 U1114 ( .A(n2271), .B(n2279), .C(n1587), .Y(n1218) );
  OAI21X1 U1116 ( .A(n2270), .B(n2279), .C(n348), .Y(n1219) );
  OAI21X1 U1118 ( .A(n2269), .B(n2279), .C(n1249), .Y(n1220) );
  OAI21X1 U1120 ( .A(n2268), .B(n2279), .C(n43), .Y(n1221) );
  OAI21X1 U1122 ( .A(n2267), .B(n2279), .C(n88), .Y(n1222) );
  OAI21X1 U1124 ( .A(n2266), .B(n2279), .C(n1470), .Y(n1223) );
  OAI21X1 U1126 ( .A(n2265), .B(n2279), .C(n1506), .Y(n1224) );
  OAI21X1 U1128 ( .A(n2264), .B(n2279), .C(n1337), .Y(n1225) );
  OAI21X1 U1130 ( .A(n2263), .B(n2279), .C(n1369), .Y(n1226) );
  NOR3X1 U1133 ( .A(n2345), .B(n2344), .C(n2346), .Y(n244) );
  NOR3X1 U1134 ( .A(n2347), .B(n658), .C(n2348), .Y(n536) );
  OAI21X1 U1135 ( .A(n2348), .B(n1711), .C(n1545), .Y(n1227) );
  OAI21X1 U1137 ( .A(n2347), .B(n1711), .C(n1505), .Y(n1228) );
  OAI21X1 U1139 ( .A(n2346), .B(n1711), .C(n1469), .Y(n1229) );
  OAI21X1 U1141 ( .A(n2345), .B(n1711), .C(n1435), .Y(n1230) );
  OAI21X1 U1143 ( .A(n2344), .B(n1711), .C(n1401), .Y(n1231) );
  AOI22X1 U1147 ( .A(n58), .B(n2262), .C(n23), .D(n667), .Y(n665) );
  AOI22X1 U1148 ( .A(n57), .B(n2262), .C(n22), .D(n667), .Y(n668) );
  AOI22X1 U1149 ( .A(n56), .B(n2262), .C(n21), .D(n667), .Y(n669) );
  AOI22X1 U1150 ( .A(n55), .B(n2262), .C(n20), .D(n667), .Y(n670) );
  AOI22X1 U1151 ( .A(n2240), .B(n2262), .C(n2311), .D(n667), .Y(n671) );
  AOI22X1 U1152 ( .A(data_out[15]), .B(n2261), .C(n24), .D(n2262), .Y(n672) );
  AOI22X1 U1153 ( .A(data_out[14]), .B(n2261), .C(n25), .D(n2262), .Y(n673) );
  AOI22X1 U1154 ( .A(data_out[13]), .B(n2261), .C(n26), .D(n2262), .Y(n674) );
  AOI22X1 U1155 ( .A(data_out[12]), .B(n2261), .C(n27), .D(n2262), .Y(n675) );
  AOI22X1 U1156 ( .A(data_out[11]), .B(n2261), .C(n28), .D(n2262), .Y(n676) );
  AOI22X1 U1157 ( .A(data_out[10]), .B(n2261), .C(n29), .D(n2262), .Y(n677) );
  AOI22X1 U1158 ( .A(data_out[9]), .B(n2261), .C(n30), .D(n2262), .Y(n678) );
  AOI22X1 U1159 ( .A(data_out[8]), .B(n2261), .C(n31), .D(n2262), .Y(n679) );
  AOI22X1 U1160 ( .A(data_out[7]), .B(n2261), .C(n32), .D(n1583), .Y(n680) );
  AOI22X1 U1161 ( .A(data_out[6]), .B(n2261), .C(n33), .D(n2262), .Y(n681) );
  AOI22X1 U1162 ( .A(data_out[5]), .B(n2261), .C(n34), .D(n1583), .Y(n682) );
  AOI22X1 U1163 ( .A(data_out[4]), .B(n2261), .C(n35), .D(n2262), .Y(n683) );
  AOI22X1 U1164 ( .A(data_out[3]), .B(n2261), .C(n36), .D(n2262), .Y(n684) );
  AOI22X1 U1165 ( .A(data_out[2]), .B(n2261), .C(n37), .D(n2262), .Y(n685) );
  AOI22X1 U1166 ( .A(data_out[1]), .B(n2261), .C(n38), .D(n2262), .Y(n686) );
  AOI22X1 U1167 ( .A(data_out[0]), .B(n2261), .C(n39), .D(n2262), .Y(n687) );
  OAI21X1 U1169 ( .A(n690), .B(n2349), .C(n1436), .Y(n1232) );
  AOI22X1 U1170 ( .A(n81), .B(n692), .C(n69), .D(n693), .Y(n691) );
  OAI21X1 U1171 ( .A(n690), .B(n2317), .C(n1540), .Y(n1233) );
  AOI22X1 U1172 ( .A(n80), .B(n692), .C(n68), .D(n693), .Y(n694) );
  OAI21X1 U1173 ( .A(n690), .B(n2318), .C(n1504), .Y(n1234) );
  AOI22X1 U1174 ( .A(n79), .B(n692), .C(n67), .D(n693), .Y(n695) );
  OAI21X1 U1175 ( .A(n690), .B(n2350), .C(n1582), .Y(n1235) );
  AOI22X1 U1176 ( .A(n78), .B(n692), .C(n66), .D(n693), .Y(n696) );
  OAI21X1 U1177 ( .A(n690), .B(n77), .C(n1402), .Y(n1236) );
  AOI22X1 U1178 ( .A(n77), .B(n692), .C(n77), .D(n693), .Y(n697) );
  OAI21X1 U1179 ( .A(n1585), .B(n2343), .C(n1584), .Y(n1237) );
  NAND3X1 U1181 ( .A(n1586), .B(n2312), .C(n1625), .Y(n698) );
  NAND3X1 U1182 ( .A(n702), .B(n2319), .C(n703), .Y(n701) );
  NOR3X1 U1183 ( .A(n1707), .B(fillcount[3]), .C(fillcount[2]), .Y(n703) );
  OAI21X1 U1185 ( .A(n690), .B(n2342), .C(n1623), .Y(n1238) );
  AOI22X1 U1186 ( .A(n82), .B(n692), .C(n70), .D(n693), .Y(n705) );
  OAI21X1 U1188 ( .A(n1543), .B(n2341), .C(n1542), .Y(n1239) );
  NAND3X1 U1190 ( .A(n1544), .B(n2312), .C(n1710), .Y(n708) );
  NAND3X1 U1191 ( .A(get), .B(n2343), .C(n707), .Y(n688) );
  NAND3X1 U1192 ( .A(n1624), .B(n663), .C(n713), .Y(n710) );
  NOR3X1 U1193 ( .A(n1664), .B(fillcount[5]), .C(n2349), .Y(n713) );
  NAND3X1 U1196 ( .A(n711), .B(n2343), .C(get), .Y(n689) );
  HAX1 add_45_U1_1_1 ( .A(fillcount[1]), .B(fillcount[0]), .YC(add_45_carry[2]), .YS(n66) );
  HAX1 add_45_U1_1_2 ( .A(fillcount[2]), .B(add_45_carry[2]), .YC(
        add_45_carry[3]), .YS(n67) );
  HAX1 add_45_U1_1_3 ( .A(fillcount[3]), .B(add_45_carry[3]), .YC(
        add_45_carry[4]), .YS(n68) );
  HAX1 add_45_U1_1_4 ( .A(fillcount[4]), .B(add_45_carry[4]), .YC(
        add_45_carry[5]), .YS(n69) );
  HAX1 r308_U1_1_1 ( .A(n20), .B(n2311), .YC(r308_carry[2]), .YS(n55) );
  HAX1 r308_U1_1_2 ( .A(n21), .B(r308_carry[2]), .YC(r308_carry[3]), .YS(n56)
         );
  HAX1 r308_U1_1_3 ( .A(n22), .B(r308_carry[3]), .YC(r308_carry[4]), .YS(n57)
         );
  HAX1 r307_U1_1_1 ( .A(wr_ptr[1]), .B(wr_ptr[0]), .YC(r307_carry[2]), .YS(n50) );
  HAX1 r307_U1_1_2 ( .A(wr_ptr[2]), .B(r307_carry[2]), .YC(r307_carry[3]), 
        .YS(n51) );
  HAX1 r307_U1_1_3 ( .A(wr_ptr[3]), .B(r307_carry[3]), .YC(r307_carry[4]), 
        .YS(n52) );
  OR2X1 U3 ( .A(n1541), .B(reset), .Y(n664) );
  OR2X1 U4 ( .A(n1667), .B(n663), .Y(n690) );
  OR2X1 U5 ( .A(n1709), .B(fillcount[4]), .Y(n2316) );
  AND2X1 U6 ( .A(n1585), .B(n1667), .Y(n699) );
  AND2X1 U7 ( .A(n663), .B(n1543), .Y(n709) );
  AND2X1 U8 ( .A(n1625), .B(n664), .Y(n658) );
  AND2X1 U9 ( .A(n706), .B(n1541), .Y(n663) );
  AND2X1 U10 ( .A(put), .B(n2341), .Y(n711) );
  BUFX2 U11 ( .A(n687), .Y(n1) );
  BUFX2 U12 ( .A(n686), .Y(n2) );
  BUFX2 U13 ( .A(n685), .Y(n3) );
  BUFX2 U14 ( .A(n684), .Y(n4) );
  BUFX2 U15 ( .A(n683), .Y(n5) );
  BUFX2 U16 ( .A(n682), .Y(n6) );
  BUFX2 U17 ( .A(n681), .Y(n7) );
  BUFX2 U18 ( .A(n680), .Y(n8) );
  BUFX2 U19 ( .A(n679), .Y(n9) );
  BUFX2 U20 ( .A(n678), .Y(n10) );
  BUFX2 U21 ( .A(n677), .Y(n11) );
  BUFX2 U22 ( .A(n676), .Y(n12) );
  BUFX2 U23 ( .A(n675), .Y(n13) );
  BUFX2 U24 ( .A(n674), .Y(n14) );
  BUFX2 U25 ( .A(n673), .Y(n15) );
  BUFX2 U26 ( .A(n672), .Y(n16) );
  BUFX2 U27 ( .A(n671), .Y(n17) );
  BUFX2 U28 ( .A(n670), .Y(n18) );
  BUFX2 U29 ( .A(n669), .Y(n40) );
  BUFX2 U30 ( .A(n668), .Y(n41) );
  BUFX2 U31 ( .A(n665), .Y(n42) );
  AND2X1 U32 ( .A(fifo_array[506]), .B(n2279), .Y(n650) );
  INVX1 U33 ( .A(n650), .Y(n43) );
  AND2X1 U34 ( .A(fifo_array[491]), .B(n2280), .Y(n634) );
  INVX1 U35 ( .A(n634), .Y(n44) );
  AND2X1 U36 ( .A(fifo_array[478]), .B(n2281), .Y(n620) );
  INVX1 U37 ( .A(n620), .Y(n45) );
  AND2X1 U38 ( .A(fifo_array[463]), .B(n2282), .Y(n604) );
  INVX1 U39 ( .A(n604), .Y(n46) );
  AND2X1 U40 ( .A(fifo_array[403]), .B(n2285), .Y(n541) );
  INVX1 U41 ( .A(n541), .Y(n47) );
  AND2X1 U42 ( .A(fifo_array[388]), .B(n2286), .Y(n524) );
  INVX1 U43 ( .A(n524), .Y(n48) );
  AND2X1 U44 ( .A(fifo_array[373]), .B(n2287), .Y(n508) );
  INVX1 U45 ( .A(n508), .Y(n49) );
  AND2X1 U46 ( .A(fifo_array[358]), .B(n2288), .Y(n492) );
  INVX1 U47 ( .A(n492), .Y(n54) );
  AND2X1 U48 ( .A(fifo_array[343]), .B(n2289), .Y(n476) );
  INVX1 U49 ( .A(n476), .Y(n59) );
  AND2X1 U50 ( .A(fifo_array[328]), .B(n2290), .Y(n460) );
  INVX1 U51 ( .A(n460), .Y(n60) );
  AND2X1 U52 ( .A(fifo_array[313]), .B(n2291), .Y(n444) );
  INVX1 U53 ( .A(n444), .Y(n61) );
  AND2X1 U54 ( .A(fifo_array[298]), .B(n2292), .Y(n428) );
  INVX1 U55 ( .A(n428), .Y(n62) );
  AND2X1 U56 ( .A(fifo_array[283]), .B(n2293), .Y(n412) );
  INVX1 U57 ( .A(n412), .Y(n63) );
  AND2X1 U58 ( .A(fifo_array[270]), .B(n2294), .Y(n397) );
  INVX1 U59 ( .A(n397), .Y(n64) );
  AND2X1 U60 ( .A(fifo_array[255]), .B(n2295), .Y(n381) );
  INVX1 U61 ( .A(n381), .Y(n65) );
  AND2X1 U62 ( .A(fifo_array[195]), .B(n2298), .Y(n318) );
  INVX1 U63 ( .A(n318), .Y(n71) );
  AND2X1 U64 ( .A(fifo_array[180]), .B(n2299), .Y(n302) );
  INVX1 U65 ( .A(n302), .Y(n72) );
  AND2X1 U66 ( .A(fifo_array[165]), .B(n2300), .Y(n286) );
  INVX1 U68 ( .A(n286), .Y(n73) );
  AND2X1 U70 ( .A(fifo_array[150]), .B(n2301), .Y(n270) );
  INVX1 U72 ( .A(n270), .Y(n74) );
  AND2X1 U74 ( .A(fifo_array[135]), .B(n2302), .Y(n253) );
  INVX1 U76 ( .A(n253), .Y(n75) );
  AND2X1 U78 ( .A(fifo_array[120]), .B(n2303), .Y(n236) );
  INVX1 U80 ( .A(n236), .Y(n76) );
  AND2X1 U82 ( .A(fifo_array[105]), .B(n2304), .Y(n219) );
  INVX1 U84 ( .A(n219), .Y(n83) );
  AND2X1 U86 ( .A(fifo_array[90]), .B(n2305), .Y(n202) );
  INVX1 U88 ( .A(n202), .Y(n84) );
  AND2X1 U90 ( .A(fifo_array[75]), .B(n2306), .Y(n185) );
  INVX1 U92 ( .A(n185), .Y(n85) );
  AND2X1 U94 ( .A(fifo_array[62]), .B(n2307), .Y(n170) );
  INVX1 U96 ( .A(n170), .Y(n86) );
  AND2X1 U98 ( .A(fifo_array[47]), .B(n2308), .Y(n153) );
  INVX1 U99 ( .A(n153), .Y(n87) );
  AND2X1 U101 ( .A(fifo_array[507]), .B(n2279), .Y(n651) );
  INVX1 U103 ( .A(n651), .Y(n88) );
  AND2X1 U105 ( .A(fifo_array[490]), .B(n2280), .Y(n633) );
  INVX1 U107 ( .A(n633), .Y(n89) );
  AND2X1 U109 ( .A(fifo_array[479]), .B(n2281), .Y(n621) );
  INVX1 U111 ( .A(n621), .Y(n90) );
  AND2X1 U113 ( .A(fifo_array[462]), .B(n2282), .Y(n603) );
  INVX1 U115 ( .A(n603), .Y(n91) );
  AND2X1 U117 ( .A(fifo_array[402]), .B(n2285), .Y(n540) );
  INVX1 U119 ( .A(n540), .Y(n92) );
  AND2X1 U121 ( .A(fifo_array[389]), .B(n2286), .Y(n525) );
  INVX1 U123 ( .A(n525), .Y(n93) );
  AND2X1 U125 ( .A(fifo_array[372]), .B(n2287), .Y(n507) );
  INVX1 U127 ( .A(n507), .Y(n94) );
  AND2X1 U129 ( .A(fifo_array[359]), .B(n2288), .Y(n493) );
  INVX1 U131 ( .A(n493), .Y(n95) );
  AND2X1 U132 ( .A(fifo_array[342]), .B(n2289), .Y(n475) );
  INVX1 U134 ( .A(n475), .Y(n96) );
  AND2X1 U136 ( .A(fifo_array[329]), .B(n2290), .Y(n461) );
  INVX1 U138 ( .A(n461), .Y(n97) );
  AND2X1 U140 ( .A(fifo_array[312]), .B(n2291), .Y(n443) );
  INVX1 U142 ( .A(n443), .Y(n98) );
  AND2X1 U144 ( .A(fifo_array[299]), .B(n2292), .Y(n429) );
  INVX1 U146 ( .A(n429), .Y(n99) );
  AND2X1 U148 ( .A(fifo_array[282]), .B(n2293), .Y(n411) );
  INVX1 U150 ( .A(n411), .Y(n100) );
  AND2X1 U152 ( .A(fifo_array[271]), .B(n2294), .Y(n398) );
  INVX1 U154 ( .A(n398), .Y(n119) );
  AND2X1 U156 ( .A(fifo_array[254]), .B(n2295), .Y(n380) );
  INVX1 U158 ( .A(n380), .Y(n137) );
  AND2X1 U160 ( .A(fifo_array[194]), .B(n2298), .Y(n317) );
  INVX1 U162 ( .A(n317), .Y(n155) );
  AND2X1 U164 ( .A(fifo_array[181]), .B(n2299), .Y(n303) );
  INVX1 U165 ( .A(n303), .Y(n173) );
  AND2X1 U167 ( .A(fifo_array[164]), .B(n2300), .Y(n285) );
  INVX1 U169 ( .A(n285), .Y(n191) );
  AND2X1 U171 ( .A(fifo_array[151]), .B(n2301), .Y(n271) );
  INVX1 U173 ( .A(n271), .Y(n209) );
  AND2X1 U175 ( .A(fifo_array[134]), .B(n2302), .Y(n252) );
  INVX1 U177 ( .A(n252), .Y(n227) );
  AND2X1 U179 ( .A(fifo_array[121]), .B(n2303), .Y(n237) );
  INVX1 U181 ( .A(n237), .Y(n245) );
  AND2X1 U183 ( .A(fifo_array[104]), .B(n2304), .Y(n218) );
  INVX1 U185 ( .A(n218), .Y(n263) );
  AND2X1 U187 ( .A(fifo_array[91]), .B(n2305), .Y(n203) );
  INVX1 U189 ( .A(n203), .Y(n280) );
  AND2X1 U191 ( .A(fifo_array[74]), .B(n2306), .Y(n184) );
  INVX1 U193 ( .A(n184), .Y(n297) );
  AND2X1 U195 ( .A(fifo_array[63]), .B(n2307), .Y(n171) );
  INVX1 U197 ( .A(n171), .Y(n314) );
  AND2X1 U198 ( .A(fifo_array[46]), .B(n2308), .Y(n152) );
  INVX1 U200 ( .A(n152), .Y(n331) );
  AND2X1 U202 ( .A(fifo_array[504]), .B(n2279), .Y(n648) );
  INVX1 U204 ( .A(n648), .Y(n348) );
  AND2X1 U206 ( .A(fifo_array[489]), .B(n2280), .Y(n632) );
  INVX1 U208 ( .A(n632), .Y(n365) );
  AND2X1 U210 ( .A(fifo_array[446]), .B(n2283), .Y(n586) );
  INVX1 U212 ( .A(n586), .Y(n382) );
  AND2X1 U214 ( .A(fifo_array[431]), .B(n2284), .Y(n570) );
  INVX1 U216 ( .A(n570), .Y(n400) );
  AND2X1 U218 ( .A(fifo_array[413]), .B(n2285), .Y(n551) );
  INVX1 U220 ( .A(n551), .Y(n417) );
  AND2X1 U222 ( .A(fifo_array[401]), .B(n2285), .Y(n539) );
  INVX1 U224 ( .A(n539), .Y(n434) );
  AND2X1 U226 ( .A(fifo_array[390]), .B(n2286), .Y(n526) );
  INVX1 U228 ( .A(n526), .Y(n451) );
  AND2X1 U230 ( .A(fifo_array[375]), .B(n2287), .Y(n510) );
  INVX1 U231 ( .A(n510), .Y(n468) );
  AND2X1 U233 ( .A(fifo_array[356]), .B(n2288), .Y(n490) );
  INVX1 U235 ( .A(n490), .Y(n485) );
  AND2X1 U237 ( .A(fifo_array[341]), .B(n2289), .Y(n474) );
  INVX1 U239 ( .A(n474), .Y(n502) );
  AND2X1 U241 ( .A(fifo_array[330]), .B(n2290), .Y(n462) );
  INVX1 U243 ( .A(n462), .Y(n519) );
  AND2X1 U245 ( .A(fifo_array[315]), .B(n2291), .Y(n446) );
  INVX1 U247 ( .A(n446), .Y(n537) );
  AND2X1 U249 ( .A(fifo_array[296]), .B(n2292), .Y(n426) );
  INVX1 U251 ( .A(n426), .Y(n554) );
  AND2X1 U253 ( .A(fifo_array[281]), .B(n2293), .Y(n410) );
  INVX1 U255 ( .A(n410), .Y(n571) );
  AND2X1 U257 ( .A(fifo_array[238]), .B(n2296), .Y(n363) );
  INVX1 U259 ( .A(n363), .Y(n588) );
  AND2X1 U261 ( .A(fifo_array[223]), .B(n2297), .Y(n347) );
  INVX1 U263 ( .A(n347), .Y(n605) );
  AND2X1 U264 ( .A(fifo_array[205]), .B(n2298), .Y(n328) );
  INVX1 U266 ( .A(n328), .Y(n622) );
  AND2X1 U268 ( .A(fifo_array[193]), .B(n2298), .Y(n316) );
  INVX1 U270 ( .A(n316), .Y(n639) );
  AND2X1 U272 ( .A(fifo_array[182]), .B(n2299), .Y(n304) );
  INVX1 U274 ( .A(n304), .Y(n666) );
  AND2X1 U276 ( .A(fifo_array[167]), .B(n2300), .Y(n288) );
  INVX1 U278 ( .A(n288), .Y(n1240) );
  AND2X1 U280 ( .A(fifo_array[148]), .B(n2301), .Y(n268) );
  INVX1 U282 ( .A(n268), .Y(n1241) );
  AND2X1 U284 ( .A(fifo_array[133]), .B(n2302), .Y(n251) );
  INVX1 U286 ( .A(n251), .Y(n1242) );
  AND2X1 U288 ( .A(fifo_array[122]), .B(n2303), .Y(n238) );
  INVX1 U290 ( .A(n238), .Y(n1243) );
  AND2X1 U292 ( .A(fifo_array[107]), .B(n2304), .Y(n221) );
  INVX1 U294 ( .A(n221), .Y(n1244) );
  AND2X1 U296 ( .A(fifo_array[88]), .B(n2305), .Y(n200) );
  INVX1 U297 ( .A(n200), .Y(n1245) );
  AND2X1 U299 ( .A(fifo_array[73]), .B(n2306), .Y(n183) );
  INVX1 U301 ( .A(n183), .Y(n1246) );
  AND2X1 U303 ( .A(fifo_array[30]), .B(n2309), .Y(n134) );
  INVX1 U305 ( .A(n134), .Y(n1247) );
  AND2X1 U307 ( .A(fifo_array[15]), .B(n2310), .Y(n116) );
  INVX1 U309 ( .A(n116), .Y(n1248) );
  AND2X1 U311 ( .A(fifo_array[505]), .B(n2279), .Y(n649) );
  INVX1 U313 ( .A(n649), .Y(n1249) );
  AND2X1 U315 ( .A(fifo_array[488]), .B(n2280), .Y(n631) );
  INVX1 U317 ( .A(n631), .Y(n1250) );
  AND2X1 U319 ( .A(fifo_array[447]), .B(n2283), .Y(n587) );
  INVX1 U321 ( .A(n587), .Y(n1251) );
  AND2X1 U323 ( .A(fifo_array[430]), .B(n2284), .Y(n569) );
  INVX1 U325 ( .A(n569), .Y(n1252) );
  AND2X1 U327 ( .A(fifo_array[412]), .B(n2285), .Y(n550) );
  INVX1 U329 ( .A(n550), .Y(n1253) );
  AND2X1 U330 ( .A(fifo_array[400]), .B(n2285), .Y(n538) );
  INVX1 U333 ( .A(n538), .Y(n1254) );
  AND2X1 U335 ( .A(fifo_array[391]), .B(n2286), .Y(n527) );
  INVX1 U337 ( .A(n527), .Y(n1255) );
  AND2X1 U339 ( .A(fifo_array[374]), .B(n2287), .Y(n509) );
  INVX1 U341 ( .A(n509), .Y(n1256) );
  AND2X1 U343 ( .A(fifo_array[357]), .B(n2288), .Y(n491) );
  INVX1 U345 ( .A(n491), .Y(n1257) );
  AND2X1 U347 ( .A(fifo_array[340]), .B(n2289), .Y(n473) );
  INVX1 U349 ( .A(n473), .Y(n1258) );
  AND2X1 U351 ( .A(fifo_array[331]), .B(n2290), .Y(n463) );
  INVX1 U353 ( .A(n463), .Y(n1259) );
  AND2X1 U355 ( .A(fifo_array[314]), .B(n2291), .Y(n445) );
  INVX1 U357 ( .A(n445), .Y(n1260) );
  AND2X1 U359 ( .A(fifo_array[297]), .B(n2292), .Y(n427) );
  INVX1 U361 ( .A(n427), .Y(n1261) );
  AND2X1 U363 ( .A(fifo_array[280]), .B(n2293), .Y(n409) );
  INVX1 U364 ( .A(n409), .Y(n1262) );
  AND2X1 U366 ( .A(fifo_array[239]), .B(n2296), .Y(n364) );
  INVX1 U368 ( .A(n364), .Y(n1263) );
  AND2X1 U370 ( .A(fifo_array[222]), .B(n2297), .Y(n346) );
  INVX1 U372 ( .A(n346), .Y(n1264) );
  AND2X1 U374 ( .A(fifo_array[204]), .B(n2298), .Y(n327) );
  INVX1 U376 ( .A(n327), .Y(n1265) );
  AND2X1 U378 ( .A(fifo_array[192]), .B(n2298), .Y(n315) );
  INVX1 U380 ( .A(n315), .Y(n1266) );
  AND2X1 U382 ( .A(fifo_array[183]), .B(n2299), .Y(n305) );
  INVX1 U384 ( .A(n305), .Y(n1267) );
  AND2X1 U386 ( .A(fifo_array[166]), .B(n2300), .Y(n287) );
  INVX1 U388 ( .A(n287), .Y(n1268) );
  AND2X1 U390 ( .A(fifo_array[149]), .B(n2301), .Y(n269) );
  INVX1 U392 ( .A(n269), .Y(n1269) );
  AND2X1 U394 ( .A(fifo_array[132]), .B(n2302), .Y(n250) );
  INVX1 U396 ( .A(n250), .Y(n1270) );
  AND2X1 U397 ( .A(fifo_array[123]), .B(n2303), .Y(n239) );
  INVX1 U399 ( .A(n239), .Y(n1271) );
  AND2X1 U401 ( .A(fifo_array[106]), .B(n2304), .Y(n220) );
  INVX1 U403 ( .A(n220), .Y(n1272) );
  AND2X1 U405 ( .A(fifo_array[89]), .B(n2305), .Y(n201) );
  INVX1 U407 ( .A(n201), .Y(n1273) );
  AND2X1 U409 ( .A(fifo_array[72]), .B(n2306), .Y(n182) );
  INVX1 U411 ( .A(n182), .Y(n1274) );
  AND2X1 U413 ( .A(fifo_array[31]), .B(n2309), .Y(n135) );
  INVX1 U415 ( .A(n135), .Y(n1275) );
  AND2X1 U417 ( .A(fifo_array[14]), .B(n2310), .Y(n115) );
  INVX1 U419 ( .A(n115), .Y(n1276) );
  AND2X1 U421 ( .A(fifo_array[472]), .B(n2281), .Y(n614) );
  INVX1 U423 ( .A(n614), .Y(n1277) );
  AND2X1 U425 ( .A(fifo_array[457]), .B(n2282), .Y(n598) );
  INVX1 U427 ( .A(n598), .Y(n1278) );
  AND2X1 U429 ( .A(fifo_array[442]), .B(n2283), .Y(n582) );
  INVX1 U430 ( .A(n582), .Y(n1279) );
  AND2X1 U432 ( .A(fifo_array[427]), .B(n2284), .Y(n566) );
  INVX1 U434 ( .A(n566), .Y(n1280) );
  AND2X1 U436 ( .A(fifo_array[407]), .B(n2285), .Y(n545) );
  INVX1 U438 ( .A(n545), .Y(n1281) );
  AND2X1 U440 ( .A(fifo_array[396]), .B(n2286), .Y(n532) );
  INVX1 U442 ( .A(n532), .Y(n1282) );
  AND2X1 U444 ( .A(fifo_array[384]), .B(n2286), .Y(n520) );
  INVX1 U446 ( .A(n520), .Y(n1283) );
  AND2X1 U448 ( .A(fifo_array[381]), .B(n2287), .Y(n516) );
  INVX1 U450 ( .A(n516), .Y(n1284) );
  AND2X1 U452 ( .A(fifo_array[369]), .B(n2287), .Y(n504) );
  INVX1 U454 ( .A(n504), .Y(n1285) );
  AND2X1 U456 ( .A(fifo_array[354]), .B(n2288), .Y(n488) );
  INVX1 U458 ( .A(n488), .Y(n1286) );
  AND2X1 U460 ( .A(fifo_array[339]), .B(n2289), .Y(n472) );
  INVX1 U462 ( .A(n472), .Y(n1287) );
  AND2X1 U463 ( .A(fifo_array[334]), .B(n2290), .Y(n466) );
  INVX1 U465 ( .A(n466), .Y(n1288) );
  AND2X1 U467 ( .A(fifo_array[319]), .B(n2291), .Y(n450) );
  INVX1 U469 ( .A(n450), .Y(n1289) );
  AND2X1 U471 ( .A(fifo_array[264]), .B(n2294), .Y(n391) );
  INVX1 U473 ( .A(n391), .Y(n1290) );
  AND2X1 U475 ( .A(fifo_array[249]), .B(n2295), .Y(n375) );
  INVX1 U477 ( .A(n375), .Y(n1291) );
  AND2X1 U479 ( .A(fifo_array[234]), .B(n2296), .Y(n359) );
  INVX1 U481 ( .A(n359), .Y(n1292) );
  AND2X1 U483 ( .A(fifo_array[219]), .B(n2297), .Y(n343) );
  INVX1 U485 ( .A(n343), .Y(n1293) );
  AND2X1 U487 ( .A(fifo_array[199]), .B(n2298), .Y(n322) );
  INVX1 U489 ( .A(n322), .Y(n1294) );
  AND2X1 U491 ( .A(fifo_array[188]), .B(n2299), .Y(n310) );
  INVX1 U493 ( .A(n310), .Y(n1295) );
  AND2X1 U495 ( .A(fifo_array[176]), .B(n2299), .Y(n298) );
  INVX1 U496 ( .A(n298), .Y(n1296) );
  AND2X1 U498 ( .A(fifo_array[173]), .B(n2300), .Y(n294) );
  INVX1 U500 ( .A(n294), .Y(n1297) );
  AND2X1 U502 ( .A(fifo_array[161]), .B(n2300), .Y(n282) );
  INVX1 U504 ( .A(n282), .Y(n1298) );
  AND2X1 U506 ( .A(fifo_array[146]), .B(n2301), .Y(n266) );
  INVX1 U508 ( .A(n266), .Y(n1299) );
  AND2X1 U510 ( .A(fifo_array[131]), .B(n2302), .Y(n249) );
  INVX1 U512 ( .A(n249), .Y(n1300) );
  AND2X1 U514 ( .A(fifo_array[126]), .B(n2303), .Y(n242) );
  INVX1 U516 ( .A(n242), .Y(n1301) );
  AND2X1 U518 ( .A(fifo_array[111]), .B(n2304), .Y(n225) );
  INVX1 U520 ( .A(n225), .Y(n1302) );
  AND2X1 U522 ( .A(fifo_array[56]), .B(n2307), .Y(n164) );
  INVX1 U524 ( .A(n164), .Y(n1303) );
  AND2X1 U526 ( .A(fifo_array[41]), .B(n2308), .Y(n147) );
  INVX1 U528 ( .A(n147), .Y(n1304) );
  AND2X1 U529 ( .A(fifo_array[26]), .B(n2309), .Y(n130) );
  INVX1 U531 ( .A(n130), .Y(n1305) );
  AND2X1 U533 ( .A(fifo_array[11]), .B(n2310), .Y(n112) );
  INVX1 U535 ( .A(n112), .Y(n1306) );
  AND2X1 U537 ( .A(fifo_array[473]), .B(n2281), .Y(n615) );
  INVX1 U539 ( .A(n615), .Y(n1307) );
  AND2X1 U541 ( .A(fifo_array[456]), .B(n2282), .Y(n597) );
  INVX1 U543 ( .A(n597), .Y(n1308) );
  AND2X1 U545 ( .A(fifo_array[443]), .B(n2283), .Y(n583) );
  INVX1 U547 ( .A(n583), .Y(n1309) );
  AND2X1 U549 ( .A(fifo_array[426]), .B(n2284), .Y(n565) );
  INVX1 U551 ( .A(n565), .Y(n1310) );
  AND2X1 U553 ( .A(fifo_array[406]), .B(n2285), .Y(n544) );
  INVX1 U555 ( .A(n544), .Y(n1311) );
  AND2X1 U557 ( .A(fifo_array[397]), .B(n2286), .Y(n533) );
  INVX1 U559 ( .A(n533), .Y(n1312) );
  AND2X1 U561 ( .A(fifo_array[385]), .B(n2286), .Y(n521) );
  INVX1 U562 ( .A(n521), .Y(n1313) );
  AND2X1 U564 ( .A(fifo_array[380]), .B(n2287), .Y(n515) );
  INVX1 U566 ( .A(n515), .Y(n1314) );
  AND2X1 U568 ( .A(fifo_array[368]), .B(n2287), .Y(n503) );
  INVX1 U570 ( .A(n503), .Y(n1315) );
  AND2X1 U572 ( .A(fifo_array[355]), .B(n2288), .Y(n489) );
  INVX1 U574 ( .A(n489), .Y(n1316) );
  AND2X1 U576 ( .A(fifo_array[338]), .B(n2289), .Y(n471) );
  INVX1 U578 ( .A(n471), .Y(n1317) );
  AND2X1 U580 ( .A(fifo_array[335]), .B(n2290), .Y(n467) );
  INVX1 U582 ( .A(n467), .Y(n1318) );
  AND2X1 U584 ( .A(fifo_array[318]), .B(n2291), .Y(n449) );
  INVX1 U586 ( .A(n449), .Y(n1319) );
  AND2X1 U588 ( .A(fifo_array[265]), .B(n2294), .Y(n392) );
  INVX1 U590 ( .A(n392), .Y(n1320) );
  AND2X1 U592 ( .A(fifo_array[248]), .B(n2295), .Y(n374) );
  INVX1 U594 ( .A(n374), .Y(n1321) );
  AND2X1 U595 ( .A(fifo_array[235]), .B(n2296), .Y(n360) );
  INVX1 U598 ( .A(n360), .Y(n1322) );
  AND2X1 U600 ( .A(fifo_array[218]), .B(n2297), .Y(n342) );
  INVX1 U602 ( .A(n342), .Y(n1323) );
  AND2X1 U604 ( .A(fifo_array[198]), .B(n2298), .Y(n321) );
  INVX1 U606 ( .A(n321), .Y(n1324) );
  AND2X1 U608 ( .A(fifo_array[189]), .B(n2299), .Y(n311) );
  INVX1 U610 ( .A(n311), .Y(n1325) );
  AND2X1 U612 ( .A(fifo_array[177]), .B(n2299), .Y(n299) );
  INVX1 U614 ( .A(n299), .Y(n1326) );
  AND2X1 U616 ( .A(fifo_array[172]), .B(n2300), .Y(n293) );
  INVX1 U618 ( .A(n293), .Y(n1327) );
  AND2X1 U620 ( .A(fifo_array[160]), .B(n2300), .Y(n281) );
  INVX1 U622 ( .A(n281), .Y(n1328) );
  AND2X1 U624 ( .A(fifo_array[147]), .B(n2301), .Y(n267) );
  INVX1 U626 ( .A(n267), .Y(n1329) );
  AND2X1 U628 ( .A(fifo_array[130]), .B(n2302), .Y(n248) );
  INVX1 U629 ( .A(n248), .Y(n1330) );
  AND2X1 U631 ( .A(fifo_array[127]), .B(n2303), .Y(n243) );
  INVX1 U633 ( .A(n243), .Y(n1331) );
  AND2X1 U635 ( .A(fifo_array[110]), .B(n2304), .Y(n224) );
  INVX1 U637 ( .A(n224), .Y(n1332) );
  AND2X1 U639 ( .A(fifo_array[57]), .B(n2307), .Y(n165) );
  INVX1 U641 ( .A(n165), .Y(n1333) );
  AND2X1 U643 ( .A(fifo_array[40]), .B(n2308), .Y(n146) );
  INVX1 U645 ( .A(n146), .Y(n1334) );
  AND2X1 U647 ( .A(fifo_array[27]), .B(n2309), .Y(n131) );
  INVX1 U649 ( .A(n131), .Y(n1335) );
  AND2X1 U651 ( .A(fifo_array[10]), .B(n2310), .Y(n111) );
  INVX1 U653 ( .A(n111), .Y(n1336) );
  AND2X1 U655 ( .A(fifo_array[510]), .B(n2279), .Y(n654) );
  INVX1 U657 ( .A(n654), .Y(n1337) );
  AND2X1 U659 ( .A(fifo_array[495]), .B(n2280), .Y(n638) );
  INVX1 U661 ( .A(n638), .Y(n1338) );
  AND2X1 U662 ( .A(fifo_array[474]), .B(n2281), .Y(n616) );
  INVX1 U664 ( .A(n616), .Y(n1339) );
  AND2X1 U666 ( .A(fifo_array[459]), .B(n2282), .Y(n600) );
  INVX1 U668 ( .A(n600), .Y(n1340) );
  AND2X1 U670 ( .A(fifo_array[440]), .B(n2283), .Y(n580) );
  INVX1 U672 ( .A(n580), .Y(n1341) );
  AND2X1 U674 ( .A(fifo_array[425]), .B(n2284), .Y(n564) );
  INVX1 U676 ( .A(n564), .Y(n1342) );
  AND2X1 U678 ( .A(fifo_array[405]), .B(n2285), .Y(n543) );
  INVX1 U680 ( .A(n543), .Y(n1343) );
  AND2X1 U682 ( .A(fifo_array[386]), .B(n2286), .Y(n522) );
  INVX1 U684 ( .A(n522), .Y(n1344) );
  AND2X1 U686 ( .A(fifo_array[371]), .B(n2287), .Y(n506) );
  INVX1 U688 ( .A(n506), .Y(n1345) );
  AND2X1 U690 ( .A(fifo_array[364]), .B(n2288), .Y(n498) );
  INVX1 U692 ( .A(n498), .Y(n1346) );
  AND2X1 U694 ( .A(fifo_array[352]), .B(n2288), .Y(n486) );
  INVX1 U695 ( .A(n486), .Y(n1347) );
  AND2X1 U697 ( .A(fifo_array[349]), .B(n2289), .Y(n482) );
  INVX1 U699 ( .A(n482), .Y(n1348) );
  AND2X1 U701 ( .A(fifo_array[337]), .B(n2289), .Y(n470) );
  INVX1 U703 ( .A(n470), .Y(n1349) );
  AND2X1 U705 ( .A(fifo_array[302]), .B(n2292), .Y(n432) );
  INVX1 U707 ( .A(n432), .Y(n1350) );
  AND2X1 U709 ( .A(fifo_array[287]), .B(n2293), .Y(n416) );
  INVX1 U711 ( .A(n416), .Y(n1351) );
  AND2X1 U713 ( .A(fifo_array[266]), .B(n2294), .Y(n393) );
  INVX1 U715 ( .A(n393), .Y(n1352) );
  AND2X1 U717 ( .A(fifo_array[251]), .B(n2295), .Y(n377) );
  INVX1 U719 ( .A(n377), .Y(n1353) );
  AND2X1 U721 ( .A(fifo_array[232]), .B(n2296), .Y(n357) );
  INVX1 U723 ( .A(n357), .Y(n1354) );
  AND2X1 U725 ( .A(fifo_array[217]), .B(n2297), .Y(n341) );
  INVX1 U727 ( .A(n341), .Y(n1355) );
  AND2X1 U728 ( .A(fifo_array[197]), .B(n2298), .Y(n320) );
  INVX1 U730 ( .A(n320), .Y(n1356) );
  AND2X1 U732 ( .A(fifo_array[178]), .B(n2299), .Y(n300) );
  INVX1 U734 ( .A(n300), .Y(n1357) );
  AND2X1 U736 ( .A(fifo_array[163]), .B(n2300), .Y(n284) );
  INVX1 U738 ( .A(n284), .Y(n1358) );
  AND2X1 U740 ( .A(fifo_array[156]), .B(n2301), .Y(n276) );
  INVX1 U742 ( .A(n276), .Y(n1359) );
  AND2X1 U744 ( .A(fifo_array[144]), .B(n2301), .Y(n264) );
  INVX1 U746 ( .A(n264), .Y(n1360) );
  AND2X1 U748 ( .A(fifo_array[141]), .B(n2302), .Y(n259) );
  INVX1 U750 ( .A(n259), .Y(n1361) );
  AND2X1 U752 ( .A(fifo_array[129]), .B(n2302), .Y(n247) );
  INVX1 U754 ( .A(n247), .Y(n1362) );
  AND2X1 U756 ( .A(fifo_array[94]), .B(n2305), .Y(n206) );
  INVX1 U758 ( .A(n206), .Y(n1363) );
  AND2X1 U760 ( .A(fifo_array[79]), .B(n2306), .Y(n189) );
  INVX1 U761 ( .A(n189), .Y(n1364) );
  AND2X1 U763 ( .A(fifo_array[58]), .B(n2307), .Y(n166) );
  INVX1 U765 ( .A(n166), .Y(n1365) );
  AND2X1 U767 ( .A(fifo_array[43]), .B(n2308), .Y(n149) );
  INVX1 U769 ( .A(n149), .Y(n1366) );
  AND2X1 U771 ( .A(fifo_array[24]), .B(n2309), .Y(n128) );
  INVX1 U773 ( .A(n128), .Y(n1367) );
  AND2X1 U775 ( .A(fifo_array[9]), .B(n2310), .Y(n110) );
  INVX1 U777 ( .A(n110), .Y(n1368) );
  AND2X1 U779 ( .A(fifo_array[511]), .B(n2279), .Y(n655) );
  INVX1 U781 ( .A(n655), .Y(n1369) );
  AND2X1 U783 ( .A(fifo_array[494]), .B(n2280), .Y(n637) );
  INVX1 U785 ( .A(n637), .Y(n1370) );
  AND2X1 U787 ( .A(fifo_array[475]), .B(n2281), .Y(n617) );
  INVX1 U789 ( .A(n617), .Y(n1371) );
  AND2X1 U791 ( .A(fifo_array[458]), .B(n2282), .Y(n599) );
  INVX1 U793 ( .A(n599), .Y(n1372) );
  AND2X1 U794 ( .A(fifo_array[441]), .B(n2283), .Y(n581) );
  INVX1 U796 ( .A(n581), .Y(n1373) );
  AND2X1 U798 ( .A(fifo_array[424]), .B(n2284), .Y(n563) );
  INVX1 U800 ( .A(n563), .Y(n1374) );
  AND2X1 U802 ( .A(fifo_array[404]), .B(n2285), .Y(n542) );
  INVX1 U804 ( .A(n542), .Y(n1375) );
  AND2X1 U806 ( .A(fifo_array[387]), .B(n2286), .Y(n523) );
  INVX1 U808 ( .A(n523), .Y(n1376) );
  AND2X1 U810 ( .A(fifo_array[370]), .B(n2287), .Y(n505) );
  INVX1 U812 ( .A(n505), .Y(n1377) );
  AND2X1 U814 ( .A(fifo_array[365]), .B(n2288), .Y(n499) );
  INVX1 U816 ( .A(n499), .Y(n1378) );
  AND2X1 U818 ( .A(fifo_array[353]), .B(n2288), .Y(n487) );
  INVX1 U820 ( .A(n487), .Y(n1379) );
  AND2X1 U822 ( .A(fifo_array[348]), .B(n2289), .Y(n481) );
  INVX1 U824 ( .A(n481), .Y(n1380) );
  AND2X1 U826 ( .A(fifo_array[336]), .B(n2289), .Y(n469) );
  INVX1 U827 ( .A(n469), .Y(n1381) );
  AND2X1 U829 ( .A(fifo_array[303]), .B(n2292), .Y(n433) );
  INVX1 U831 ( .A(n433), .Y(n1382) );
  AND2X1 U833 ( .A(fifo_array[286]), .B(n2293), .Y(n415) );
  INVX1 U835 ( .A(n415), .Y(n1383) );
  AND2X1 U837 ( .A(fifo_array[267]), .B(n2294), .Y(n394) );
  INVX1 U839 ( .A(n394), .Y(n1384) );
  AND2X1 U841 ( .A(fifo_array[250]), .B(n2295), .Y(n376) );
  INVX1 U843 ( .A(n376), .Y(n1385) );
  AND2X1 U845 ( .A(fifo_array[233]), .B(n2296), .Y(n358) );
  INVX1 U847 ( .A(n358), .Y(n1386) );
  AND2X1 U849 ( .A(fifo_array[216]), .B(n2297), .Y(n340) );
  INVX1 U851 ( .A(n340), .Y(n1387) );
  AND2X1 U853 ( .A(fifo_array[196]), .B(n2298), .Y(n319) );
  INVX1 U855 ( .A(n319), .Y(n1388) );
  AND2X1 U857 ( .A(fifo_array[179]), .B(n2299), .Y(n301) );
  INVX1 U859 ( .A(n301), .Y(n1389) );
  AND2X1 U860 ( .A(fifo_array[162]), .B(n2300), .Y(n283) );
  INVX1 U863 ( .A(n283), .Y(n1390) );
  AND2X1 U865 ( .A(fifo_array[157]), .B(n2301), .Y(n277) );
  INVX1 U867 ( .A(n277), .Y(n1391) );
  AND2X1 U869 ( .A(fifo_array[145]), .B(n2301), .Y(n265) );
  INVX1 U871 ( .A(n265), .Y(n1392) );
  AND2X1 U873 ( .A(fifo_array[140]), .B(n2302), .Y(n258) );
  INVX1 U875 ( .A(n258), .Y(n1393) );
  AND2X1 U877 ( .A(fifo_array[128]), .B(n2302), .Y(n246) );
  INVX1 U879 ( .A(n246), .Y(n1394) );
  AND2X1 U881 ( .A(fifo_array[95]), .B(n2305), .Y(n207) );
  INVX1 U883 ( .A(n207), .Y(n1395) );
  AND2X1 U885 ( .A(fifo_array[78]), .B(n2306), .Y(n188) );
  INVX1 U887 ( .A(n188), .Y(n1396) );
  AND2X1 U889 ( .A(fifo_array[59]), .B(n2307), .Y(n167) );
  INVX1 U891 ( .A(n167), .Y(n1397) );
  AND2X1 U893 ( .A(fifo_array[42]), .B(n2308), .Y(n148) );
  INVX1 U894 ( .A(n148), .Y(n1398) );
  AND2X1 U897 ( .A(fifo_array[25]), .B(n2309), .Y(n129) );
  INVX1 U899 ( .A(n129), .Y(n1399) );
  AND2X1 U901 ( .A(fifo_array[8]), .B(n2310), .Y(n109) );
  INVX1 U903 ( .A(n109), .Y(n1400) );
  AND2X1 U905 ( .A(n2344), .B(n1668), .Y(n662) );
  INVX1 U907 ( .A(n662), .Y(n1401) );
  BUFX2 U909 ( .A(n697), .Y(n1402) );
  AND2X1 U911 ( .A(fifo_array[498]), .B(n2279), .Y(n642) );
  INVX1 U913 ( .A(n642), .Y(n1403) );
  AND2X1 U915 ( .A(fifo_array[483]), .B(n2280), .Y(n626) );
  INVX1 U917 ( .A(n626), .Y(n1404) );
  AND2X1 U919 ( .A(fifo_array[468]), .B(n2281), .Y(n610) );
  INVX1 U921 ( .A(n610), .Y(n1405) );
  AND2X1 U923 ( .A(fifo_array[453]), .B(n2282), .Y(n594) );
  INVX1 U925 ( .A(n594), .Y(n1406) );
  AND2X1 U927 ( .A(fifo_array[438]), .B(n2283), .Y(n578) );
  INVX1 U928 ( .A(n578), .Y(n1407) );
  AND2X1 U931 ( .A(fifo_array[423]), .B(n2284), .Y(n562) );
  INVX1 U933 ( .A(n562), .Y(n1408) );
  AND2X1 U935 ( .A(fifo_array[411]), .B(n2285), .Y(n549) );
  INVX1 U937 ( .A(n549), .Y(n1409) );
  AND2X1 U939 ( .A(fifo_array[398]), .B(n2286), .Y(n534) );
  INVX1 U941 ( .A(n534), .Y(n1410) );
  AND2X1 U943 ( .A(fifo_array[383]), .B(n2287), .Y(n518) );
  INVX1 U945 ( .A(n518), .Y(n1411) );
  AND2X1 U947 ( .A(fifo_array[332]), .B(n2290), .Y(n464) );
  INVX1 U949 ( .A(n464), .Y(n1412) );
  AND2X1 U951 ( .A(fifo_array[320]), .B(n2290), .Y(n452) );
  INVX1 U953 ( .A(n452), .Y(n1413) );
  AND2X1 U955 ( .A(fifo_array[317]), .B(n2291), .Y(n448) );
  INVX1 U957 ( .A(n448), .Y(n1414) );
  AND2X1 U959 ( .A(fifo_array[305]), .B(n2291), .Y(n436) );
  INVX1 U961 ( .A(n436), .Y(n1415) );
  AND2X1 U962 ( .A(fifo_array[290]), .B(n2292), .Y(n420) );
  INVX1 U965 ( .A(n420), .Y(n1416) );
  AND2X1 U967 ( .A(fifo_array[275]), .B(n2293), .Y(n404) );
  INVX1 U969 ( .A(n404), .Y(n1417) );
  AND2X1 U971 ( .A(fifo_array[260]), .B(n2294), .Y(n387) );
  INVX1 U973 ( .A(n387), .Y(n1418) );
  AND2X1 U975 ( .A(fifo_array[245]), .B(n2295), .Y(n371) );
  INVX1 U977 ( .A(n371), .Y(n1419) );
  AND2X1 U979 ( .A(fifo_array[230]), .B(n2296), .Y(n355) );
  INVX1 U981 ( .A(n355), .Y(n1420) );
  AND2X1 U983 ( .A(fifo_array[215]), .B(n2297), .Y(n339) );
  INVX1 U985 ( .A(n339), .Y(n1421) );
  AND2X1 U987 ( .A(fifo_array[203]), .B(n2298), .Y(n326) );
  INVX1 U989 ( .A(n326), .Y(n1422) );
  AND2X1 U991 ( .A(fifo_array[190]), .B(n2299), .Y(n312) );
  INVX1 U993 ( .A(n312), .Y(n1423) );
  AND2X1 U995 ( .A(fifo_array[175]), .B(n2300), .Y(n296) );
  INVX1 U996 ( .A(n296), .Y(n1424) );
  AND2X1 U999 ( .A(fifo_array[124]), .B(n2303), .Y(n240) );
  INVX1 U1001 ( .A(n240), .Y(n1425) );
  AND2X1 U1003 ( .A(fifo_array[112]), .B(n2303), .Y(n228) );
  INVX1 U1005 ( .A(n228), .Y(n1426) );
  AND2X1 U1007 ( .A(fifo_array[109]), .B(n2304), .Y(n223) );
  INVX1 U1009 ( .A(n223), .Y(n1427) );
  AND2X1 U1011 ( .A(fifo_array[97]), .B(n2304), .Y(n211) );
  INVX1 U1013 ( .A(n211), .Y(n1428) );
  AND2X1 U1015 ( .A(fifo_array[82]), .B(n2305), .Y(n194) );
  INVX1 U1017 ( .A(n194), .Y(n1429) );
  AND2X1 U1019 ( .A(fifo_array[67]), .B(n2306), .Y(n177) );
  INVX1 U1021 ( .A(n177), .Y(n1430) );
  AND2X1 U1023 ( .A(fifo_array[52]), .B(n2307), .Y(n160) );
  INVX1 U1025 ( .A(n160), .Y(n1431) );
  AND2X1 U1027 ( .A(fifo_array[37]), .B(n2308), .Y(n143) );
  INVX1 U1029 ( .A(n143), .Y(n1432) );
  AND2X1 U1030 ( .A(fifo_array[22]), .B(n2309), .Y(n126) );
  INVX1 U1033 ( .A(n126), .Y(n1433) );
  AND2X1 U1035 ( .A(fifo_array[7]), .B(n2310), .Y(n108) );
  INVX1 U1037 ( .A(n108), .Y(n1434) );
  AND2X1 U1039 ( .A(n50), .B(n1668), .Y(n661) );
  INVX1 U1041 ( .A(n661), .Y(n1435) );
  BUFX2 U1043 ( .A(n691), .Y(n1436) );
  AND2X1 U1045 ( .A(fifo_array[499]), .B(n2279), .Y(n643) );
  INVX1 U1047 ( .A(n643), .Y(n1437) );
  AND2X1 U1049 ( .A(fifo_array[482]), .B(n2280), .Y(n625) );
  INVX1 U1051 ( .A(n625), .Y(n1438) );
  AND2X1 U1053 ( .A(fifo_array[469]), .B(n2281), .Y(n611) );
  INVX1 U1055 ( .A(n611), .Y(n1439) );
  AND2X1 U1057 ( .A(fifo_array[452]), .B(n2282), .Y(n593) );
  INVX1 U1059 ( .A(n593), .Y(n1440) );
  AND2X1 U1061 ( .A(fifo_array[439]), .B(n2283), .Y(n579) );
  INVX1 U1063 ( .A(n579), .Y(n1441) );
  AND2X1 U1064 ( .A(fifo_array[422]), .B(n2284), .Y(n561) );
  INVX1 U1067 ( .A(n561), .Y(n1442) );
  AND2X1 U1069 ( .A(fifo_array[410]), .B(n2285), .Y(n548) );
  INVX1 U1071 ( .A(n548), .Y(n1443) );
  AND2X1 U1073 ( .A(fifo_array[399]), .B(n2286), .Y(n535) );
  INVX1 U1075 ( .A(n535), .Y(n1444) );
  AND2X1 U1077 ( .A(fifo_array[382]), .B(n2287), .Y(n517) );
  INVX1 U1079 ( .A(n517), .Y(n1445) );
  AND2X1 U1081 ( .A(fifo_array[333]), .B(n2290), .Y(n465) );
  INVX1 U1083 ( .A(n465), .Y(n1446) );
  AND2X1 U1085 ( .A(fifo_array[321]), .B(n2290), .Y(n453) );
  INVX1 U1087 ( .A(n453), .Y(n1447) );
  AND2X1 U1089 ( .A(fifo_array[316]), .B(n2291), .Y(n447) );
  INVX1 U1091 ( .A(n447), .Y(n1448) );
  AND2X1 U1093 ( .A(fifo_array[304]), .B(n2291), .Y(n435) );
  INVX1 U1095 ( .A(n435), .Y(n1449) );
  AND2X1 U1097 ( .A(fifo_array[291]), .B(n2292), .Y(n421) );
  INVX1 U1098 ( .A(n421), .Y(n1450) );
  AND2X1 U1101 ( .A(fifo_array[274]), .B(n2293), .Y(n403) );
  INVX1 U1103 ( .A(n403), .Y(n1451) );
  AND2X1 U1105 ( .A(fifo_array[261]), .B(n2294), .Y(n388) );
  INVX1 U1107 ( .A(n388), .Y(n1452) );
  AND2X1 U1109 ( .A(fifo_array[244]), .B(n2295), .Y(n370) );
  INVX1 U1111 ( .A(n370), .Y(n1453) );
  AND2X1 U1113 ( .A(fifo_array[231]), .B(n2296), .Y(n356) );
  INVX1 U1115 ( .A(n356), .Y(n1454) );
  AND2X1 U1117 ( .A(fifo_array[214]), .B(n2297), .Y(n338) );
  INVX1 U1119 ( .A(n338), .Y(n1455) );
  AND2X1 U1121 ( .A(fifo_array[202]), .B(n2298), .Y(n325) );
  INVX1 U1123 ( .A(n325), .Y(n1456) );
  AND2X1 U1125 ( .A(fifo_array[191]), .B(n2299), .Y(n313) );
  INVX1 U1127 ( .A(n313), .Y(n1457) );
  AND2X1 U1129 ( .A(fifo_array[174]), .B(n2300), .Y(n295) );
  INVX1 U1131 ( .A(n295), .Y(n1458) );
  AND2X1 U1132 ( .A(fifo_array[125]), .B(n2303), .Y(n241) );
  INVX1 U1136 ( .A(n241), .Y(n1459) );
  AND2X1 U1138 ( .A(fifo_array[113]), .B(n2303), .Y(n229) );
  INVX1 U1140 ( .A(n229), .Y(n1460) );
  AND2X1 U1142 ( .A(fifo_array[108]), .B(n2304), .Y(n222) );
  INVX1 U1144 ( .A(n222), .Y(n1461) );
  AND2X1 U1145 ( .A(fifo_array[96]), .B(n2304), .Y(n210) );
  INVX1 U1146 ( .A(n210), .Y(n1462) );
  AND2X1 U1168 ( .A(fifo_array[83]), .B(n2305), .Y(n195) );
  INVX1 U1180 ( .A(n195), .Y(n1463) );
  AND2X1 U1184 ( .A(fifo_array[66]), .B(n2306), .Y(n176) );
  INVX1 U1187 ( .A(n176), .Y(n1464) );
  AND2X1 U1189 ( .A(fifo_array[53]), .B(n2307), .Y(n161) );
  INVX1 U1194 ( .A(n161), .Y(n1465) );
  AND2X1 U1195 ( .A(fifo_array[36]), .B(n2308), .Y(n142) );
  INVX1 U1197 ( .A(n142), .Y(n1466) );
  AND2X1 U1198 ( .A(fifo_array[23]), .B(n2309), .Y(n127) );
  INVX1 U1199 ( .A(n127), .Y(n1467) );
  AND2X1 U1200 ( .A(fifo_array[6]), .B(n2310), .Y(n107) );
  INVX1 U1201 ( .A(n107), .Y(n1468) );
  AND2X1 U1202 ( .A(n1665), .B(n2312), .Y(n707) );
  AND2X1 U1203 ( .A(n51), .B(n1668), .Y(n660) );
  INVX1 U1204 ( .A(n660), .Y(n1469) );
  AND2X1 U1205 ( .A(fifo_array[508]), .B(n2279), .Y(n652) );
  INVX1 U1206 ( .A(n652), .Y(n1470) );
  AND2X1 U1207 ( .A(fifo_array[496]), .B(n2279), .Y(n640) );
  INVX1 U1208 ( .A(n640), .Y(n1471) );
  AND2X1 U1209 ( .A(fifo_array[493]), .B(n2280), .Y(n636) );
  INVX1 U1210 ( .A(n636), .Y(n1472) );
  AND2X1 U1211 ( .A(fifo_array[481]), .B(n2280), .Y(n624) );
  INVX1 U1212 ( .A(n624), .Y(n1473) );
  AND2X1 U1213 ( .A(fifo_array[470]), .B(n2281), .Y(n612) );
  INVX1 U1214 ( .A(n612), .Y(n1474) );
  AND2X1 U1215 ( .A(fifo_array[455]), .B(n2282), .Y(n596) );
  INVX1 U1216 ( .A(n596), .Y(n1475) );
  AND2X1 U1217 ( .A(fifo_array[436]), .B(n2283), .Y(n576) );
  INVX1 U1218 ( .A(n576), .Y(n1476) );
  AND2X1 U1219 ( .A(fifo_array[421]), .B(n2284), .Y(n560) );
  INVX1 U1220 ( .A(n560), .Y(n1477) );
  AND2X1 U1221 ( .A(fifo_array[409]), .B(n2285), .Y(n547) );
  INVX1 U1222 ( .A(n547), .Y(n1478) );
  AND2X1 U1223 ( .A(fifo_array[366]), .B(n2288), .Y(n500) );
  INVX1 U1224 ( .A(n500), .Y(n1479) );
  AND2X1 U1225 ( .A(fifo_array[351]), .B(n2289), .Y(n484) );
  INVX1 U1226 ( .A(n484), .Y(n1480) );
  AND2X1 U1227 ( .A(fifo_array[322]), .B(n2290), .Y(n454) );
  INVX1 U1228 ( .A(n454), .Y(n1481) );
  AND2X1 U1229 ( .A(fifo_array[307]), .B(n2291), .Y(n438) );
  INVX1 U1230 ( .A(n438), .Y(n1482) );
  AND2X1 U1231 ( .A(fifo_array[300]), .B(n2292), .Y(n430) );
  INVX1 U1232 ( .A(n430), .Y(n1483) );
  AND2X1 U1233 ( .A(fifo_array[288]), .B(n2292), .Y(n418) );
  INVX1 U1234 ( .A(n418), .Y(n1484) );
  AND2X1 U1235 ( .A(fifo_array[285]), .B(n2293), .Y(n414) );
  INVX1 U1236 ( .A(n414), .Y(n1485) );
  AND2X1 U1237 ( .A(fifo_array[273]), .B(n2293), .Y(n402) );
  INVX1 U1238 ( .A(n402), .Y(n1486) );
  AND2X1 U1239 ( .A(fifo_array[262]), .B(n2294), .Y(n389) );
  INVX1 U1240 ( .A(n389), .Y(n1487) );
  AND2X1 U1241 ( .A(fifo_array[247]), .B(n2295), .Y(n373) );
  INVX1 U1242 ( .A(n373), .Y(n1488) );
  AND2X1 U1243 ( .A(fifo_array[228]), .B(n2296), .Y(n353) );
  INVX1 U1244 ( .A(n353), .Y(n1489) );
  AND2X1 U1245 ( .A(fifo_array[213]), .B(n2297), .Y(n337) );
  INVX1 U1246 ( .A(n337), .Y(n1490) );
  AND2X1 U1247 ( .A(fifo_array[201]), .B(n2298), .Y(n324) );
  INVX1 U1248 ( .A(n324), .Y(n1491) );
  AND2X1 U1249 ( .A(fifo_array[158]), .B(n2301), .Y(n278) );
  INVX1 U1250 ( .A(n278), .Y(n1492) );
  AND2X1 U1251 ( .A(fifo_array[143]), .B(n2302), .Y(n261) );
  INVX1 U1252 ( .A(n261), .Y(n1493) );
  AND2X1 U1253 ( .A(fifo_array[114]), .B(n2303), .Y(n230) );
  INVX1 U1254 ( .A(n230), .Y(n1494) );
  AND2X1 U1255 ( .A(fifo_array[99]), .B(n2304), .Y(n213) );
  INVX1 U1256 ( .A(n213), .Y(n1495) );
  AND2X1 U1257 ( .A(fifo_array[92]), .B(n2305), .Y(n204) );
  INVX1 U1258 ( .A(n204), .Y(n1496) );
  AND2X1 U1259 ( .A(fifo_array[80]), .B(n2305), .Y(n192) );
  INVX1 U1260 ( .A(n192), .Y(n1497) );
  AND2X1 U1261 ( .A(fifo_array[77]), .B(n2306), .Y(n187) );
  INVX1 U1262 ( .A(n187), .Y(n1498) );
  AND2X1 U1263 ( .A(fifo_array[65]), .B(n2306), .Y(n175) );
  INVX1 U1264 ( .A(n175), .Y(n1499) );
  AND2X1 U1265 ( .A(fifo_array[54]), .B(n2307), .Y(n162) );
  INVX1 U1266 ( .A(n162), .Y(n1500) );
  AND2X1 U1267 ( .A(fifo_array[39]), .B(n2308), .Y(n145) );
  INVX1 U1268 ( .A(n145), .Y(n1501) );
  AND2X1 U1269 ( .A(fifo_array[20]), .B(n2309), .Y(n124) );
  INVX1 U1270 ( .A(n124), .Y(n1502) );
  AND2X1 U1271 ( .A(fifo_array[5]), .B(n2310), .Y(n106) );
  INVX1 U1272 ( .A(n106), .Y(n1503) );
  BUFX2 U1273 ( .A(n695), .Y(n1504) );
  AND2X1 U1274 ( .A(n52), .B(n1668), .Y(n659) );
  INVX1 U1275 ( .A(n659), .Y(n1505) );
  AND2X1 U1276 ( .A(fifo_array[509]), .B(n2279), .Y(n653) );
  INVX1 U1277 ( .A(n653), .Y(n1506) );
  AND2X1 U1278 ( .A(fifo_array[497]), .B(n2279), .Y(n641) );
  INVX1 U1279 ( .A(n641), .Y(n1507) );
  AND2X1 U1280 ( .A(fifo_array[492]), .B(n2280), .Y(n635) );
  INVX1 U1281 ( .A(n635), .Y(n1508) );
  AND2X1 U1282 ( .A(fifo_array[480]), .B(n2280), .Y(n623) );
  INVX1 U1283 ( .A(n623), .Y(n1509) );
  AND2X1 U1284 ( .A(fifo_array[471]), .B(n2281), .Y(n613) );
  INVX1 U1285 ( .A(n613), .Y(n1510) );
  AND2X1 U1286 ( .A(fifo_array[454]), .B(n2282), .Y(n595) );
  INVX1 U1287 ( .A(n595), .Y(n1511) );
  AND2X1 U1288 ( .A(fifo_array[437]), .B(n2283), .Y(n577) );
  INVX1 U1289 ( .A(n577), .Y(n1512) );
  AND2X1 U1290 ( .A(fifo_array[420]), .B(n2284), .Y(n559) );
  INVX1 U1291 ( .A(n559), .Y(n1513) );
  AND2X1 U1292 ( .A(fifo_array[408]), .B(n2285), .Y(n546) );
  INVX1 U1293 ( .A(n546), .Y(n1514) );
  AND2X1 U1294 ( .A(fifo_array[367]), .B(n2288), .Y(n501) );
  INVX1 U1295 ( .A(n501), .Y(n1515) );
  AND2X1 U1296 ( .A(fifo_array[350]), .B(n2289), .Y(n483) );
  INVX1 U1297 ( .A(n483), .Y(n1516) );
  AND2X1 U1298 ( .A(fifo_array[323]), .B(n2290), .Y(n455) );
  INVX1 U1299 ( .A(n455), .Y(n1517) );
  AND2X1 U1300 ( .A(fifo_array[306]), .B(n2291), .Y(n437) );
  INVX1 U1301 ( .A(n437), .Y(n1518) );
  AND2X1 U1302 ( .A(fifo_array[301]), .B(n2292), .Y(n431) );
  INVX1 U1303 ( .A(n431), .Y(n1519) );
  AND2X1 U1304 ( .A(fifo_array[289]), .B(n2292), .Y(n419) );
  INVX1 U1305 ( .A(n419), .Y(n1520) );
  AND2X1 U1306 ( .A(fifo_array[284]), .B(n2293), .Y(n413) );
  INVX1 U1307 ( .A(n413), .Y(n1521) );
  AND2X1 U1308 ( .A(fifo_array[272]), .B(n2293), .Y(n401) );
  INVX1 U1309 ( .A(n401), .Y(n1522) );
  AND2X1 U1310 ( .A(fifo_array[263]), .B(n2294), .Y(n390) );
  INVX1 U1311 ( .A(n390), .Y(n1523) );
  AND2X1 U1312 ( .A(fifo_array[246]), .B(n2295), .Y(n372) );
  INVX1 U1313 ( .A(n372), .Y(n1524) );
  AND2X1 U1314 ( .A(fifo_array[229]), .B(n2296), .Y(n354) );
  INVX1 U1315 ( .A(n354), .Y(n1525) );
  AND2X1 U1316 ( .A(fifo_array[212]), .B(n2297), .Y(n336) );
  INVX1 U1317 ( .A(n336), .Y(n1526) );
  AND2X1 U1318 ( .A(fifo_array[200]), .B(n2298), .Y(n323) );
  INVX1 U1319 ( .A(n323), .Y(n1527) );
  AND2X1 U1320 ( .A(fifo_array[159]), .B(n2301), .Y(n279) );
  INVX1 U1321 ( .A(n279), .Y(n1528) );
  AND2X1 U1322 ( .A(fifo_array[142]), .B(n2302), .Y(n260) );
  INVX1 U1323 ( .A(n260), .Y(n1529) );
  AND2X1 U1324 ( .A(fifo_array[115]), .B(n2303), .Y(n231) );
  INVX1 U1325 ( .A(n231), .Y(n1530) );
  AND2X1 U1326 ( .A(fifo_array[98]), .B(n2304), .Y(n212) );
  INVX1 U1327 ( .A(n212), .Y(n1531) );
  AND2X1 U1328 ( .A(fifo_array[93]), .B(n2305), .Y(n205) );
  INVX1 U1329 ( .A(n205), .Y(n1532) );
  AND2X1 U1330 ( .A(fifo_array[81]), .B(n2305), .Y(n193) );
  INVX1 U1331 ( .A(n193), .Y(n1533) );
  AND2X1 U1332 ( .A(fifo_array[76]), .B(n2306), .Y(n186) );
  INVX1 U1333 ( .A(n186), .Y(n1534) );
  AND2X1 U1334 ( .A(fifo_array[64]), .B(n2306), .Y(n174) );
  INVX1 U1335 ( .A(n174), .Y(n1535) );
  AND2X1 U1336 ( .A(fifo_array[55]), .B(n2307), .Y(n163) );
  INVX1 U1337 ( .A(n163), .Y(n1536) );
  AND2X1 U1338 ( .A(fifo_array[38]), .B(n2308), .Y(n144) );
  INVX1 U1339 ( .A(n144), .Y(n1537) );
  AND2X1 U1340 ( .A(fifo_array[21]), .B(n2309), .Y(n125) );
  INVX1 U1341 ( .A(n125), .Y(n1538) );
  AND2X1 U1342 ( .A(fifo_array[4]), .B(n2310), .Y(n105) );
  INVX1 U1343 ( .A(n105), .Y(n1539) );
  BUFX2 U1344 ( .A(n694), .Y(n1540) );
  BUFX2 U1345 ( .A(n689), .Y(n1541) );
  INVX1 U1346 ( .A(n709), .Y(n1542) );
  BUFX2 U1347 ( .A(n708), .Y(n1543) );
  BUFX2 U1348 ( .A(n710), .Y(n1544) );
  AND2X1 U1349 ( .A(n53), .B(n1668), .Y(n657) );
  INVX1 U1350 ( .A(n657), .Y(n1545) );
  AND2X1 U1351 ( .A(fifo_array[502]), .B(n2279), .Y(n646) );
  INVX1 U1352 ( .A(n646), .Y(n1546) );
  AND2X1 U1353 ( .A(fifo_array[487]), .B(n2280), .Y(n630) );
  INVX1 U1354 ( .A(n630), .Y(n1547) );
  AND2X1 U1355 ( .A(fifo_array[476]), .B(n2281), .Y(n618) );
  INVX1 U1356 ( .A(n618), .Y(n1548) );
  AND2X1 U1357 ( .A(fifo_array[464]), .B(n2281), .Y(n606) );
  INVX1 U1358 ( .A(n606), .Y(n1549) );
  AND2X1 U1359 ( .A(fifo_array[461]), .B(n2282), .Y(n602) );
  INVX1 U1360 ( .A(n602), .Y(n1550) );
  AND2X1 U1361 ( .A(fifo_array[449]), .B(n2282), .Y(n590) );
  INVX1 U1362 ( .A(n590), .Y(n1551) );
  AND2X1 U1363 ( .A(fifo_array[434]), .B(n2283), .Y(n574) );
  INVX1 U1364 ( .A(n574), .Y(n1552) );
  AND2X1 U1365 ( .A(fifo_array[419]), .B(n2284), .Y(n558) );
  INVX1 U1366 ( .A(n558), .Y(n1553) );
  AND2X1 U1367 ( .A(fifo_array[392]), .B(n2286), .Y(n528) );
  INVX1 U1368 ( .A(n528), .Y(n1554) );
  AND2X1 U1369 ( .A(fifo_array[377]), .B(n2287), .Y(n512) );
  INVX1 U1370 ( .A(n512), .Y(n1555) );
  AND2X1 U1371 ( .A(fifo_array[362]), .B(n2288), .Y(n496) );
  INVX1 U1372 ( .A(n496), .Y(n1556) );
  AND2X1 U1373 ( .A(fifo_array[347]), .B(n2289), .Y(n480) );
  INVX1 U1374 ( .A(n480), .Y(n1557) );
  AND2X1 U1375 ( .A(fifo_array[324]), .B(n2290), .Y(n456) );
  INVX1 U1376 ( .A(n456), .Y(n1558) );
  AND2X1 U1377 ( .A(fifo_array[309]), .B(n2291), .Y(n440) );
  INVX1 U1378 ( .A(n440), .Y(n1559) );
  AND2X1 U1379 ( .A(fifo_array[294]), .B(n2292), .Y(n424) );
  INVX1 U1380 ( .A(n424), .Y(n1560) );
  AND2X1 U1381 ( .A(fifo_array[279]), .B(n2293), .Y(n408) );
  INVX1 U1382 ( .A(n408), .Y(n1561) );
  AND2X1 U1383 ( .A(fifo_array[268]), .B(n2294), .Y(n395) );
  INVX1 U1384 ( .A(n395), .Y(n1562) );
  AND2X1 U1385 ( .A(fifo_array[256]), .B(n2294), .Y(n383) );
  INVX1 U1386 ( .A(n383), .Y(n1563) );
  AND2X1 U1387 ( .A(fifo_array[253]), .B(n2295), .Y(n379) );
  INVX1 U1388 ( .A(n379), .Y(n1564) );
  AND2X1 U1389 ( .A(fifo_array[241]), .B(n2295), .Y(n367) );
  INVX1 U1390 ( .A(n367), .Y(n1565) );
  AND2X1 U1391 ( .A(fifo_array[226]), .B(n2296), .Y(n351) );
  INVX1 U1392 ( .A(n351), .Y(n1566) );
  AND2X1 U1393 ( .A(fifo_array[211]), .B(n2297), .Y(n335) );
  INVX1 U1394 ( .A(n335), .Y(n1567) );
  AND2X1 U1395 ( .A(fifo_array[184]), .B(n2299), .Y(n306) );
  INVX1 U1396 ( .A(n306), .Y(n1568) );
  AND2X1 U1397 ( .A(fifo_array[169]), .B(n2300), .Y(n290) );
  INVX1 U1398 ( .A(n290), .Y(n1569) );
  AND2X1 U1399 ( .A(fifo_array[154]), .B(n2301), .Y(n274) );
  INVX1 U1400 ( .A(n274), .Y(n1570) );
  AND2X1 U1401 ( .A(fifo_array[139]), .B(n2302), .Y(n257) );
  INVX1 U1402 ( .A(n257), .Y(n1571) );
  AND2X1 U1403 ( .A(fifo_array[116]), .B(n2303), .Y(n232) );
  INVX1 U1404 ( .A(n232), .Y(n1572) );
  AND2X1 U1405 ( .A(fifo_array[101]), .B(n2304), .Y(n215) );
  INVX1 U1406 ( .A(n215), .Y(n1573) );
  AND2X1 U1407 ( .A(fifo_array[86]), .B(n2305), .Y(n198) );
  INVX1 U1408 ( .A(n198), .Y(n1574) );
  AND2X1 U1409 ( .A(fifo_array[71]), .B(n2306), .Y(n181) );
  INVX1 U1410 ( .A(n181), .Y(n1575) );
  AND2X1 U1411 ( .A(fifo_array[60]), .B(n2307), .Y(n168) );
  INVX1 U1412 ( .A(n168), .Y(n1576) );
  AND2X1 U1413 ( .A(fifo_array[48]), .B(n2307), .Y(n156) );
  INVX1 U1414 ( .A(n156), .Y(n1577) );
  AND2X1 U1415 ( .A(fifo_array[45]), .B(n2308), .Y(n151) );
  INVX1 U1416 ( .A(n151), .Y(n1578) );
  AND2X1 U1417 ( .A(fifo_array[33]), .B(n2308), .Y(n139) );
  INVX1 U1418 ( .A(n139), .Y(n1579) );
  AND2X1 U1419 ( .A(fifo_array[18]), .B(n2309), .Y(n122) );
  INVX1 U1420 ( .A(n122), .Y(n1580) );
  AND2X1 U1421 ( .A(fifo_array[3]), .B(n2310), .Y(n104) );
  INVX1 U1422 ( .A(n104), .Y(n1581) );
  BUFX2 U1423 ( .A(n696), .Y(n1582) );
  AND2X1 U1424 ( .A(n664), .B(n1710), .Y(n2261) );
  INVX1 U1425 ( .A(n2261), .Y(n1583) );
  INVX1 U1426 ( .A(n699), .Y(n1584) );
  BUFX2 U1427 ( .A(n698), .Y(n1585) );
  BUFX2 U1428 ( .A(n701), .Y(n1586) );
  AND2X1 U1429 ( .A(fifo_array[503]), .B(n2279), .Y(n647) );
  INVX1 U1430 ( .A(n647), .Y(n1587) );
  AND2X1 U1431 ( .A(fifo_array[486]), .B(n2280), .Y(n629) );
  INVX1 U1432 ( .A(n629), .Y(n1588) );
  AND2X1 U1433 ( .A(fifo_array[477]), .B(n2281), .Y(n619) );
  INVX1 U1434 ( .A(n619), .Y(n1589) );
  AND2X1 U1435 ( .A(fifo_array[465]), .B(n2281), .Y(n607) );
  INVX1 U1436 ( .A(n607), .Y(n1590) );
  AND2X1 U1437 ( .A(fifo_array[460]), .B(n2282), .Y(n601) );
  INVX1 U1438 ( .A(n601), .Y(n1591) );
  AND2X1 U1439 ( .A(fifo_array[448]), .B(n2282), .Y(n589) );
  INVX1 U1440 ( .A(n589), .Y(n1592) );
  AND2X1 U1441 ( .A(fifo_array[435]), .B(n2283), .Y(n575) );
  INVX1 U1442 ( .A(n575), .Y(n1593) );
  AND2X1 U1443 ( .A(fifo_array[418]), .B(n2284), .Y(n557) );
  INVX1 U1444 ( .A(n557), .Y(n1594) );
  AND2X1 U1445 ( .A(fifo_array[393]), .B(n2286), .Y(n529) );
  INVX1 U1446 ( .A(n529), .Y(n1595) );
  AND2X1 U1447 ( .A(fifo_array[376]), .B(n2287), .Y(n511) );
  INVX1 U1448 ( .A(n511), .Y(n1596) );
  AND2X1 U1449 ( .A(fifo_array[363]), .B(n2288), .Y(n497) );
  INVX1 U1450 ( .A(n497), .Y(n1597) );
  AND2X1 U1451 ( .A(fifo_array[346]), .B(n2289), .Y(n479) );
  INVX1 U1452 ( .A(n479), .Y(n1598) );
  AND2X1 U1453 ( .A(fifo_array[325]), .B(n2290), .Y(n457) );
  INVX1 U1454 ( .A(n457), .Y(n1599) );
  AND2X1 U1455 ( .A(fifo_array[308]), .B(n2291), .Y(n439) );
  INVX1 U1456 ( .A(n439), .Y(n1600) );
  AND2X1 U1457 ( .A(fifo_array[295]), .B(n2292), .Y(n425) );
  INVX1 U1458 ( .A(n425), .Y(n1601) );
  AND2X1 U1459 ( .A(fifo_array[278]), .B(n2293), .Y(n407) );
  INVX1 U1460 ( .A(n407), .Y(n1602) );
  AND2X1 U1461 ( .A(fifo_array[269]), .B(n2294), .Y(n396) );
  INVX1 U1462 ( .A(n396), .Y(n1603) );
  AND2X1 U1463 ( .A(fifo_array[257]), .B(n2294), .Y(n384) );
  INVX1 U1464 ( .A(n384), .Y(n1604) );
  AND2X1 U1465 ( .A(fifo_array[252]), .B(n2295), .Y(n378) );
  INVX1 U1466 ( .A(n378), .Y(n1605) );
  AND2X1 U1467 ( .A(fifo_array[240]), .B(n2295), .Y(n366) );
  INVX1 U1468 ( .A(n366), .Y(n1606) );
  AND2X1 U1469 ( .A(fifo_array[227]), .B(n2296), .Y(n352) );
  INVX1 U1470 ( .A(n352), .Y(n1607) );
  AND2X1 U1471 ( .A(fifo_array[210]), .B(n2297), .Y(n334) );
  INVX1 U1472 ( .A(n334), .Y(n1608) );
  AND2X1 U1473 ( .A(fifo_array[185]), .B(n2299), .Y(n307) );
  INVX1 U1474 ( .A(n307), .Y(n1609) );
  AND2X1 U1475 ( .A(fifo_array[168]), .B(n2300), .Y(n289) );
  INVX1 U1476 ( .A(n289), .Y(n1610) );
  AND2X1 U1477 ( .A(fifo_array[155]), .B(n2301), .Y(n275) );
  INVX1 U1478 ( .A(n275), .Y(n1611) );
  AND2X1 U1479 ( .A(fifo_array[138]), .B(n2302), .Y(n256) );
  INVX1 U1480 ( .A(n256), .Y(n1612) );
  AND2X1 U1481 ( .A(fifo_array[117]), .B(n2303), .Y(n233) );
  INVX1 U1482 ( .A(n233), .Y(n1613) );
  AND2X1 U1483 ( .A(fifo_array[100]), .B(n2304), .Y(n214) );
  INVX1 U1484 ( .A(n214), .Y(n1614) );
  AND2X1 U1485 ( .A(fifo_array[87]), .B(n2305), .Y(n199) );
  INVX1 U1486 ( .A(n199), .Y(n1615) );
  AND2X1 U1487 ( .A(fifo_array[70]), .B(n2306), .Y(n180) );
  INVX1 U1488 ( .A(n180), .Y(n1616) );
  AND2X1 U1489 ( .A(fifo_array[61]), .B(n2307), .Y(n169) );
  INVX1 U1490 ( .A(n169), .Y(n1617) );
  AND2X1 U1491 ( .A(fifo_array[49]), .B(n2307), .Y(n157) );
  INVX1 U1492 ( .A(n157), .Y(n1618) );
  AND2X1 U1493 ( .A(fifo_array[44]), .B(n2308), .Y(n150) );
  INVX1 U1494 ( .A(n150), .Y(n1619) );
  AND2X1 U1495 ( .A(fifo_array[32]), .B(n2308), .Y(n138) );
  INVX1 U1496 ( .A(n138), .Y(n1620) );
  AND2X1 U1497 ( .A(fifo_array[19]), .B(n2309), .Y(n123) );
  INVX1 U1498 ( .A(n123), .Y(n1621) );
  AND2X1 U1499 ( .A(fifo_array[2]), .B(n2310), .Y(n103) );
  INVX1 U1500 ( .A(n103), .Y(n1622) );
  BUFX2 U1501 ( .A(n705), .Y(n1623) );
  OR2X1 U1502 ( .A(n77), .B(n2350), .Y(n712) );
  INVX1 U1503 ( .A(n712), .Y(n1624) );
  INVX1 U1504 ( .A(n663), .Y(n1625) );
  AND2X1 U1505 ( .A(fifo_array[500]), .B(n2279), .Y(n644) );
  INVX1 U1506 ( .A(n644), .Y(n1626) );
  AND2X1 U1507 ( .A(fifo_array[485]), .B(n2280), .Y(n628) );
  INVX1 U1508 ( .A(n628), .Y(n1627) );
  AND2X1 U1509 ( .A(fifo_array[466]), .B(n2281), .Y(n608) );
  INVX1 U1510 ( .A(n608), .Y(n1628) );
  AND2X1 U1511 ( .A(fifo_array[451]), .B(n2282), .Y(n592) );
  INVX1 U1512 ( .A(n592), .Y(n1629) );
  AND2X1 U1513 ( .A(fifo_array[444]), .B(n2283), .Y(n584) );
  INVX1 U1514 ( .A(n584), .Y(n1630) );
  AND2X1 U1515 ( .A(fifo_array[432]), .B(n2283), .Y(n572) );
  INVX1 U1516 ( .A(n572), .Y(n1631) );
  AND2X1 U1517 ( .A(fifo_array[429]), .B(n2284), .Y(n568) );
  INVX1 U1518 ( .A(n568), .Y(n1632) );
  AND2X1 U1519 ( .A(fifo_array[417]), .B(n2284), .Y(n556) );
  INVX1 U1520 ( .A(n556), .Y(n1633) );
  AND2X1 U1521 ( .A(fifo_array[415]), .B(n2285), .Y(n553) );
  INVX1 U1522 ( .A(n553), .Y(n1634) );
  AND2X1 U1523 ( .A(fifo_array[394]), .B(n2286), .Y(n530) );
  INVX1 U1524 ( .A(n530), .Y(n1635) );
  AND2X1 U1525 ( .A(fifo_array[379]), .B(n2287), .Y(n514) );
  INVX1 U1526 ( .A(n514), .Y(n1636) );
  AND2X1 U1527 ( .A(fifo_array[360]), .B(n2288), .Y(n494) );
  INVX1 U1528 ( .A(n494), .Y(n1637) );
  AND2X1 U1529 ( .A(fifo_array[345]), .B(n2289), .Y(n478) );
  INVX1 U1530 ( .A(n478), .Y(n1638) );
  AND2X1 U1531 ( .A(fifo_array[326]), .B(n2290), .Y(n458) );
  INVX1 U1532 ( .A(n458), .Y(n1639) );
  AND2X1 U1533 ( .A(fifo_array[311]), .B(n2291), .Y(n442) );
  INVX1 U1534 ( .A(n442), .Y(n1640) );
  AND2X1 U1535 ( .A(fifo_array[292]), .B(n2292), .Y(n422) );
  INVX1 U1536 ( .A(n422), .Y(n1641) );
  AND2X1 U1537 ( .A(fifo_array[277]), .B(n2293), .Y(n406) );
  INVX1 U1538 ( .A(n406), .Y(n1642) );
  AND2X1 U1539 ( .A(fifo_array[258]), .B(n2294), .Y(n385) );
  INVX1 U1540 ( .A(n385), .Y(n1643) );
  AND2X1 U1541 ( .A(fifo_array[243]), .B(n2295), .Y(n369) );
  INVX1 U1542 ( .A(n369), .Y(n1644) );
  AND2X1 U1543 ( .A(fifo_array[236]), .B(n2296), .Y(n361) );
  INVX1 U1544 ( .A(n361), .Y(n1645) );
  AND2X1 U1545 ( .A(fifo_array[224]), .B(n2296), .Y(n349) );
  INVX1 U1546 ( .A(n349), .Y(n1646) );
  AND2X1 U1547 ( .A(fifo_array[221]), .B(n2297), .Y(n345) );
  INVX1 U1548 ( .A(n345), .Y(n1647) );
  AND2X1 U1549 ( .A(fifo_array[209]), .B(n2297), .Y(n333) );
  INVX1 U1550 ( .A(n333), .Y(n1648) );
  AND2X1 U1551 ( .A(fifo_array[207]), .B(n2298), .Y(n330) );
  INVX1 U1552 ( .A(n330), .Y(n1649) );
  AND2X1 U1553 ( .A(fifo_array[186]), .B(n2299), .Y(n308) );
  INVX1 U1554 ( .A(n308), .Y(n1650) );
  AND2X1 U1555 ( .A(fifo_array[171]), .B(n2300), .Y(n292) );
  INVX1 U1556 ( .A(n292), .Y(n1651) );
  AND2X1 U1557 ( .A(fifo_array[152]), .B(n2301), .Y(n272) );
  INVX1 U1558 ( .A(n272), .Y(n1652) );
  AND2X1 U1559 ( .A(fifo_array[137]), .B(n2302), .Y(n255) );
  INVX1 U1560 ( .A(n255), .Y(n1653) );
  AND2X1 U1561 ( .A(fifo_array[118]), .B(n2303), .Y(n234) );
  INVX1 U1562 ( .A(n234), .Y(n1654) );
  AND2X1 U1563 ( .A(fifo_array[103]), .B(n2304), .Y(n217) );
  INVX1 U1564 ( .A(n217), .Y(n1655) );
  AND2X1 U1565 ( .A(fifo_array[84]), .B(n2305), .Y(n196) );
  INVX1 U1566 ( .A(n196), .Y(n1656) );
  AND2X1 U1567 ( .A(fifo_array[69]), .B(n2306), .Y(n179) );
  INVX1 U1568 ( .A(n179), .Y(n1657) );
  AND2X1 U1569 ( .A(fifo_array[50]), .B(n2307), .Y(n158) );
  INVX1 U1570 ( .A(n158), .Y(n1658) );
  AND2X1 U1571 ( .A(fifo_array[35]), .B(n2308), .Y(n141) );
  INVX1 U1572 ( .A(n141), .Y(n1659) );
  AND2X1 U1573 ( .A(fifo_array[28]), .B(n2309), .Y(n132) );
  INVX1 U1574 ( .A(n132), .Y(n1660) );
  AND2X1 U1575 ( .A(fifo_array[16]), .B(n2309), .Y(n120) );
  INVX1 U1576 ( .A(n120), .Y(n1661) );
  AND2X1 U1577 ( .A(fifo_array[13]), .B(n2310), .Y(n114) );
  INVX1 U1578 ( .A(n114), .Y(n1662) );
  AND2X1 U1579 ( .A(fifo_array[1]), .B(n2310), .Y(n102) );
  INVX1 U1580 ( .A(n102), .Y(n1663) );
  AND2X1 U1581 ( .A(fillcount[2]), .B(fillcount[3]), .Y(n714) );
  INVX1 U1582 ( .A(n714), .Y(n1664) );
  INVX1 U1583 ( .A(n711), .Y(n1665) );
  AND2X1 U1584 ( .A(n2313), .B(n2318), .Y(n2314) );
  INVX1 U1585 ( .A(n2314), .Y(n1666) );
  AND2X1 U1586 ( .A(n2312), .B(n1710), .Y(n700) );
  INVX1 U1587 ( .A(n700), .Y(n1667) );
  INVX1 U1588 ( .A(n658), .Y(n1668) );
  AND2X1 U1589 ( .A(fifo_array[501]), .B(n2279), .Y(n645) );
  INVX1 U1590 ( .A(n645), .Y(n1669) );
  AND2X1 U1591 ( .A(fifo_array[484]), .B(n2280), .Y(n627) );
  INVX1 U1592 ( .A(n627), .Y(n1670) );
  AND2X1 U1593 ( .A(fifo_array[467]), .B(n2281), .Y(n609) );
  INVX1 U1594 ( .A(n609), .Y(n1671) );
  AND2X1 U1595 ( .A(fifo_array[450]), .B(n2282), .Y(n591) );
  INVX1 U1596 ( .A(n591), .Y(n1672) );
  AND2X1 U1597 ( .A(fifo_array[445]), .B(n2283), .Y(n585) );
  INVX1 U1598 ( .A(n585), .Y(n1673) );
  AND2X1 U1599 ( .A(fifo_array[433]), .B(n2283), .Y(n573) );
  INVX1 U1600 ( .A(n573), .Y(n1674) );
  AND2X1 U1601 ( .A(fifo_array[428]), .B(n2284), .Y(n567) );
  INVX1 U1602 ( .A(n567), .Y(n1675) );
  AND2X1 U1603 ( .A(fifo_array[416]), .B(n2284), .Y(n555) );
  INVX1 U1604 ( .A(n555), .Y(n1676) );
  AND2X1 U1605 ( .A(fifo_array[414]), .B(n2285), .Y(n552) );
  INVX1 U1606 ( .A(n552), .Y(n1677) );
  AND2X1 U1607 ( .A(fifo_array[395]), .B(n2286), .Y(n531) );
  INVX1 U1608 ( .A(n531), .Y(n1678) );
  AND2X1 U1609 ( .A(fifo_array[378]), .B(n2287), .Y(n513) );
  INVX1 U1610 ( .A(n513), .Y(n1679) );
  AND2X1 U1611 ( .A(fifo_array[361]), .B(n2288), .Y(n495) );
  INVX1 U1612 ( .A(n495), .Y(n1680) );
  AND2X1 U1613 ( .A(fifo_array[344]), .B(n2289), .Y(n477) );
  INVX1 U1614 ( .A(n477), .Y(n1681) );
  AND2X1 U1615 ( .A(fifo_array[327]), .B(n2290), .Y(n459) );
  INVX1 U1616 ( .A(n459), .Y(n1682) );
  AND2X1 U1617 ( .A(fifo_array[310]), .B(n2291), .Y(n441) );
  INVX1 U1618 ( .A(n441), .Y(n1683) );
  AND2X1 U1619 ( .A(fifo_array[293]), .B(n2292), .Y(n423) );
  INVX1 U1620 ( .A(n423), .Y(n1684) );
  AND2X1 U1621 ( .A(fifo_array[276]), .B(n2293), .Y(n405) );
  INVX1 U1622 ( .A(n405), .Y(n1685) );
  AND2X1 U1623 ( .A(fifo_array[259]), .B(n2294), .Y(n386) );
  INVX1 U1624 ( .A(n386), .Y(n1686) );
  AND2X1 U1625 ( .A(fifo_array[242]), .B(n2295), .Y(n368) );
  INVX1 U1626 ( .A(n368), .Y(n1687) );
  AND2X1 U1627 ( .A(fifo_array[237]), .B(n2296), .Y(n362) );
  INVX1 U1628 ( .A(n362), .Y(n1688) );
  AND2X1 U1629 ( .A(fifo_array[225]), .B(n2296), .Y(n350) );
  INVX1 U1630 ( .A(n350), .Y(n1689) );
  AND2X1 U1631 ( .A(fifo_array[220]), .B(n2297), .Y(n344) );
  INVX1 U1632 ( .A(n344), .Y(n1690) );
  AND2X1 U1633 ( .A(fifo_array[208]), .B(n2297), .Y(n332) );
  INVX1 U1634 ( .A(n332), .Y(n1691) );
  AND2X1 U1635 ( .A(fifo_array[206]), .B(n2298), .Y(n329) );
  INVX1 U1636 ( .A(n329), .Y(n1692) );
  AND2X1 U1637 ( .A(fifo_array[187]), .B(n2299), .Y(n309) );
  INVX1 U1638 ( .A(n309), .Y(n1693) );
  AND2X1 U1639 ( .A(fifo_array[170]), .B(n2300), .Y(n291) );
  INVX1 U1640 ( .A(n291), .Y(n1694) );
  AND2X1 U1641 ( .A(fifo_array[153]), .B(n2301), .Y(n273) );
  INVX1 U1642 ( .A(n273), .Y(n1695) );
  AND2X1 U1643 ( .A(fifo_array[136]), .B(n2302), .Y(n254) );
  INVX1 U1644 ( .A(n254), .Y(n1696) );
  AND2X1 U1645 ( .A(fifo_array[119]), .B(n2303), .Y(n235) );
  INVX1 U1646 ( .A(n235), .Y(n1697) );
  AND2X1 U1647 ( .A(fifo_array[102]), .B(n2304), .Y(n216) );
  INVX1 U1648 ( .A(n216), .Y(n1698) );
  AND2X1 U1649 ( .A(fifo_array[85]), .B(n2305), .Y(n197) );
  INVX1 U1650 ( .A(n197), .Y(n1699) );
  AND2X1 U1651 ( .A(fifo_array[68]), .B(n2306), .Y(n178) );
  INVX1 U1652 ( .A(n178), .Y(n1700) );
  AND2X1 U1653 ( .A(fifo_array[51]), .B(n2307), .Y(n159) );
  INVX1 U1654 ( .A(n159), .Y(n1701) );
  AND2X1 U1655 ( .A(fifo_array[34]), .B(n2308), .Y(n140) );
  INVX1 U1656 ( .A(n140), .Y(n1702) );
  AND2X1 U1657 ( .A(fifo_array[29]), .B(n2309), .Y(n133) );
  INVX1 U1658 ( .A(n133), .Y(n1703) );
  AND2X1 U1659 ( .A(fifo_array[17]), .B(n2309), .Y(n121) );
  INVX1 U1660 ( .A(n121), .Y(n1704) );
  AND2X1 U1661 ( .A(fifo_array[12]), .B(n2310), .Y(n113) );
  INVX1 U1662 ( .A(n113), .Y(n1705) );
  AND2X1 U1663 ( .A(fifo_array[0]), .B(n2310), .Y(n101) );
  INVX1 U1664 ( .A(n101), .Y(n1706) );
  AND2X1 U1665 ( .A(n2349), .B(n2342), .Y(n704) );
  INVX1 U1666 ( .A(n704), .Y(n1707) );
  AND2X1 U1667 ( .A(n2350), .B(n77), .Y(n2313) );
  INVX1 U1668 ( .A(n2313), .Y(n1708) );
  AND2X1 U1669 ( .A(n2314), .B(n2317), .Y(n2315) );
  INVX1 U1670 ( .A(n2315), .Y(n1709) );
  BUFX2 U1671 ( .A(n688), .Y(n1710) );
  AND2X1 U1672 ( .A(n658), .B(n2312), .Y(n656) );
  INVX1 U1673 ( .A(n656), .Y(n1711) );
  INVX1 U1674 ( .A(n2240), .Y(n2256) );
  INVX1 U1675 ( .A(n2240), .Y(n2255) );
  INVX1 U1676 ( .A(n2240), .Y(n2254) );
  INVX1 U1677 ( .A(n2240), .Y(n2253) );
  INVX1 U1678 ( .A(n2240), .Y(n2252) );
  INVX1 U1679 ( .A(n2240), .Y(n2251) );
  INVX1 U1680 ( .A(n2240), .Y(n2250) );
  INVX1 U1681 ( .A(n2240), .Y(n2249) );
  INVX1 U1682 ( .A(n2240), .Y(n2248) );
  INVX1 U1683 ( .A(n2240), .Y(n2247) );
  INVX1 U1684 ( .A(n2240), .Y(n2246) );
  INVX1 U1685 ( .A(n2240), .Y(n2245) );
  INVX1 U1686 ( .A(n2240), .Y(n2244) );
  INVX1 U1687 ( .A(n2240), .Y(n2243) );
  INVX1 U1688 ( .A(n2240), .Y(n2242) );
  INVX1 U1689 ( .A(n2240), .Y(n2241) );
  INVX1 U1690 ( .A(n2240), .Y(n2257) );
  INVX1 U1691 ( .A(n19), .Y(n2240) );
  AND2X1 U1692 ( .A(n706), .B(n690), .Y(n693) );
  AND2X1 U1693 ( .A(n2261), .B(n2312), .Y(n667) );
  INVX1 U1694 ( .A(n1712), .Y(n2279) );
  INVX1 U1695 ( .A(n2260), .Y(n2259) );
  INVX1 U1696 ( .A(n2260), .Y(n2258) );
  AND2X1 U1697 ( .A(n707), .B(n690), .Y(n692) );
  AND2X1 U1698 ( .A(n536), .B(n244), .Y(n1712) );
  INVX1 U1699 ( .A(n1718), .Y(n2299) );
  INVX1 U1700 ( .A(n1719), .Y(n2297) );
  INVX1 U1701 ( .A(n1713), .Y(n2296) );
  INVX1 U1702 ( .A(n1714), .Y(n2295) );
  INVX1 U1703 ( .A(n1720), .Y(n2291) );
  INVX1 U1704 ( .A(n1721), .Y(n2289) );
  INVX1 U1705 ( .A(n1715), .Y(n2288) );
  INVX1 U1706 ( .A(n1716), .Y(n2287) );
  INVX1 U1707 ( .A(n1722), .Y(n2283) );
  INVX1 U1708 ( .A(n1723), .Y(n2281) );
  INVX1 U1709 ( .A(n1717), .Y(n2280) );
  INVX1 U1710 ( .A(n1724), .Y(n2302) );
  INVX1 U1711 ( .A(n1725), .Y(n2301) );
  INVX1 U1712 ( .A(n1726), .Y(n2294) );
  INVX1 U1713 ( .A(n1727), .Y(n2293) );
  INVX1 U1714 ( .A(n1728), .Y(n2286) );
  INVX1 U1715 ( .A(n1729), .Y(n2285) );
  INVX1 U1716 ( .A(n1730), .Y(n2300) );
  INVX1 U1717 ( .A(n1731), .Y(n2298) );
  INVX1 U1718 ( .A(n1732), .Y(n2292) );
  INVX1 U1719 ( .A(n1733), .Y(n2290) );
  INVX1 U1720 ( .A(n1734), .Y(n2284) );
  INVX1 U1721 ( .A(n1735), .Y(n2282) );
  INVX1 U1722 ( .A(n1737), .Y(n2309) );
  INVX1 U1723 ( .A(n1738), .Y(n2308) );
  INVX1 U1724 ( .A(n1739), .Y(n2307) );
  INVX1 U1725 ( .A(n1740), .Y(n2306) );
  INVX1 U1726 ( .A(n1741), .Y(n2305) );
  INVX1 U1727 ( .A(n1742), .Y(n2304) );
  INVX1 U1728 ( .A(n1743), .Y(n2303) );
  INVX1 U1729 ( .A(n1736), .Y(n2310) );
  AND2X1 U1730 ( .A(n711), .B(n2312), .Y(n706) );
  INVX1 U1731 ( .A(reset), .Y(n2312) );
  INVX1 U1732 ( .A(n17), .Y(n2336) );
  AND2X1 U1733 ( .A(n262), .B(n226), .Y(n1713) );
  AND2X1 U1734 ( .A(n262), .B(n244), .Y(n1714) );
  AND2X1 U1735 ( .A(n399), .B(n226), .Y(n1715) );
  AND2X1 U1736 ( .A(n399), .B(n244), .Y(n1716) );
  AND2X1 U1737 ( .A(n536), .B(n226), .Y(n1717) );
  AND2X1 U1738 ( .A(n262), .B(n172), .Y(n1718) );
  AND2X1 U1739 ( .A(n262), .B(n208), .Y(n1719) );
  AND2X1 U1740 ( .A(n399), .B(n172), .Y(n1720) );
  AND2X1 U1741 ( .A(n399), .B(n208), .Y(n1721) );
  AND2X1 U1742 ( .A(n536), .B(n172), .Y(n1722) );
  AND2X1 U1743 ( .A(n536), .B(n208), .Y(n1723) );
  AND2X1 U1744 ( .A(n262), .B(n117), .Y(n1724) );
  AND2X1 U1745 ( .A(n262), .B(n136), .Y(n1725) );
  AND2X1 U1746 ( .A(n399), .B(n117), .Y(n1726) );
  AND2X1 U1747 ( .A(n399), .B(n136), .Y(n1727) );
  AND2X1 U1748 ( .A(n536), .B(n117), .Y(n1728) );
  AND2X1 U1749 ( .A(n536), .B(n136), .Y(n1729) );
  AND2X1 U1750 ( .A(n262), .B(n154), .Y(n1730) );
  AND2X1 U1751 ( .A(n262), .B(n190), .Y(n1731) );
  AND2X1 U1752 ( .A(n399), .B(n154), .Y(n1732) );
  AND2X1 U1753 ( .A(n399), .B(n190), .Y(n1733) );
  AND2X1 U1754 ( .A(n536), .B(n154), .Y(n1734) );
  AND2X1 U1755 ( .A(n536), .B(n190), .Y(n1735) );
  AND2X1 U1756 ( .A(n117), .B(n118), .Y(n1736) );
  AND2X1 U1757 ( .A(n136), .B(n118), .Y(n1737) );
  AND2X1 U1758 ( .A(n154), .B(n118), .Y(n1738) );
  AND2X1 U1759 ( .A(n172), .B(n118), .Y(n1739) );
  AND2X1 U1760 ( .A(n190), .B(n118), .Y(n1740) );
  AND2X1 U1761 ( .A(n208), .B(n118), .Y(n1741) );
  AND2X1 U1762 ( .A(n226), .B(n118), .Y(n1742) );
  AND2X1 U1763 ( .A(n244), .B(n118), .Y(n1743) );
  INVX1 U1764 ( .A(n1710), .Y(n2319) );
  INVX1 U1765 ( .A(data_in[0]), .Y(n2278) );
  INVX1 U1766 ( .A(data_in[1]), .Y(n2277) );
  INVX1 U1767 ( .A(data_in[2]), .Y(n2276) );
  INVX1 U1768 ( .A(data_in[3]), .Y(n2275) );
  INVX1 U1769 ( .A(data_in[4]), .Y(n2274) );
  INVX1 U1770 ( .A(data_in[5]), .Y(n2273) );
  INVX1 U1771 ( .A(data_in[6]), .Y(n2272) );
  INVX1 U1772 ( .A(data_in[7]), .Y(n2271) );
  INVX1 U1773 ( .A(data_in[8]), .Y(n2270) );
  INVX1 U1774 ( .A(data_in[9]), .Y(n2269) );
  INVX1 U1775 ( .A(data_in[10]), .Y(n2268) );
  INVX1 U1776 ( .A(data_in[11]), .Y(n2267) );
  INVX1 U1777 ( .A(data_in[12]), .Y(n2266) );
  INVX1 U1778 ( .A(data_in[13]), .Y(n2265) );
  INVX1 U1779 ( .A(data_in[14]), .Y(n2264) );
  INVX1 U1780 ( .A(data_in[15]), .Y(n2263) );
  INVX1 U1781 ( .A(n2240), .Y(n2311) );
  INVX1 U1782 ( .A(n41), .Y(n2339) );
  INVX1 U1783 ( .A(n42), .Y(n2340) );
  INVX1 U1784 ( .A(n15), .Y(n2334) );
  INVX1 U1785 ( .A(n2238), .Y(n25) );
  INVX1 U1786 ( .A(n14), .Y(n2333) );
  INVX1 U1787 ( .A(n2237), .Y(n26) );
  INVX1 U1788 ( .A(n13), .Y(n2332) );
  INVX1 U1789 ( .A(n2236), .Y(n27) );
  INVX1 U1790 ( .A(n12), .Y(n2331) );
  INVX1 U1791 ( .A(n2235), .Y(n28) );
  INVX1 U1792 ( .A(n11), .Y(n2330) );
  INVX1 U1793 ( .A(n2234), .Y(n29) );
  INVX1 U1794 ( .A(n10), .Y(n2329) );
  INVX1 U1795 ( .A(n2233), .Y(n30) );
  INVX1 U1796 ( .A(n9), .Y(n2328) );
  INVX1 U1797 ( .A(n2232), .Y(n31) );
  INVX1 U1798 ( .A(n8), .Y(n2327) );
  INVX1 U1799 ( .A(n2231), .Y(n32) );
  INVX1 U1800 ( .A(n7), .Y(n2326) );
  INVX1 U1801 ( .A(n2230), .Y(n33) );
  INVX1 U1802 ( .A(n6), .Y(n2325) );
  INVX1 U1803 ( .A(n2229), .Y(n34) );
  INVX1 U1804 ( .A(n5), .Y(n2324) );
  INVX1 U1805 ( .A(n2228), .Y(n35) );
  INVX1 U1806 ( .A(n4), .Y(n2323) );
  INVX1 U1807 ( .A(n2227), .Y(n36) );
  INVX1 U1808 ( .A(n3), .Y(n2322) );
  INVX1 U1809 ( .A(n2226), .Y(n37) );
  INVX1 U1810 ( .A(n2), .Y(n2321) );
  INVX1 U1811 ( .A(n2225), .Y(n38) );
  INVX1 U1812 ( .A(n40), .Y(n2338) );
  INVX1 U1813 ( .A(n18), .Y(n2337) );
  INVX1 U1814 ( .A(n1), .Y(n2320) );
  INVX1 U1815 ( .A(n2224), .Y(n39) );
  INVX1 U1816 ( .A(n16), .Y(n2335) );
  INVX1 U1817 ( .A(n2239), .Y(n24) );
  INVX1 U1818 ( .A(full), .Y(n2341) );
  INVX1 U1819 ( .A(wr_ptr[2]), .Y(n2346) );
  INVX1 U1820 ( .A(wr_ptr[0]), .Y(n2344) );
  INVX1 U1821 ( .A(wr_ptr[1]), .Y(n2345) );
  INVX1 U1822 ( .A(wr_ptr[4]), .Y(n2348) );
  INVX1 U1823 ( .A(wr_ptr[3]), .Y(n2347) );
  INVX1 U1824 ( .A(n20), .Y(n2260) );
  INVX1 U1825 ( .A(fillcount[4]), .Y(n2349) );
  INVX1 U1826 ( .A(fillcount[0]), .Y(n77) );
  INVX1 U1827 ( .A(fillcount[5]), .Y(n2342) );
  INVX1 U1828 ( .A(fillcount[2]), .Y(n2318) );
  INVX1 U1829 ( .A(fillcount[3]), .Y(n2317) );
  INVX1 U1830 ( .A(fillcount[1]), .Y(n2350) );
  INVX1 U1831 ( .A(empty), .Y(n2343) );
  AND2X1 U1832 ( .A(n2350), .B(fillcount[0]), .Y(n702) );
  MUX2X1 U1833 ( .B(n1745), .A(n1746), .S(n20), .Y(n1744) );
  MUX2X1 U1834 ( .B(n1748), .A(n1749), .S(n20), .Y(n1747) );
  MUX2X1 U1835 ( .B(n1751), .A(n1752), .S(n20), .Y(n1750) );
  MUX2X1 U1836 ( .B(n1754), .A(n1755), .S(n20), .Y(n1753) );
  MUX2X1 U1837 ( .B(n1757), .A(n1758), .S(n22), .Y(n1756) );
  MUX2X1 U1838 ( .B(n1760), .A(n1761), .S(n20), .Y(n1759) );
  MUX2X1 U1839 ( .B(n1763), .A(n1764), .S(n20), .Y(n1762) );
  MUX2X1 U1840 ( .B(n1766), .A(n1767), .S(n20), .Y(n1765) );
  MUX2X1 U1841 ( .B(n1769), .A(n1770), .S(n20), .Y(n1768) );
  MUX2X1 U1842 ( .B(n1772), .A(n1773), .S(n22), .Y(n1771) );
  MUX2X1 U1843 ( .B(n1775), .A(n1776), .S(n2258), .Y(n1774) );
  MUX2X1 U1844 ( .B(n1778), .A(n1779), .S(n2258), .Y(n1777) );
  MUX2X1 U1845 ( .B(n1781), .A(n1782), .S(n2258), .Y(n1780) );
  MUX2X1 U1846 ( .B(n1784), .A(n1785), .S(n2258), .Y(n1783) );
  MUX2X1 U1847 ( .B(n1787), .A(n1788), .S(n22), .Y(n1786) );
  MUX2X1 U1848 ( .B(n1790), .A(n1791), .S(n2258), .Y(n1789) );
  MUX2X1 U1849 ( .B(n1793), .A(n1794), .S(n2258), .Y(n1792) );
  MUX2X1 U1850 ( .B(n1796), .A(n1797), .S(n2258), .Y(n1795) );
  MUX2X1 U1851 ( .B(n1799), .A(n1800), .S(n2258), .Y(n1798) );
  MUX2X1 U1852 ( .B(n1802), .A(n1803), .S(n22), .Y(n1801) );
  MUX2X1 U1853 ( .B(n1805), .A(n1806), .S(n2258), .Y(n1804) );
  MUX2X1 U1854 ( .B(n1808), .A(n1809), .S(n2258), .Y(n1807) );
  MUX2X1 U1855 ( .B(n1811), .A(n1812), .S(n2258), .Y(n1810) );
  MUX2X1 U1856 ( .B(n1814), .A(n1815), .S(n2258), .Y(n1813) );
  MUX2X1 U1857 ( .B(n1817), .A(n1818), .S(n22), .Y(n1816) );
  MUX2X1 U1858 ( .B(n1820), .A(n1821), .S(n2259), .Y(n1819) );
  MUX2X1 U1859 ( .B(n1823), .A(n1824), .S(n2259), .Y(n1822) );
  MUX2X1 U1860 ( .B(n1826), .A(n1827), .S(n2259), .Y(n1825) );
  MUX2X1 U1861 ( .B(n1829), .A(n1830), .S(n2259), .Y(n1828) );
  MUX2X1 U1862 ( .B(n1832), .A(n1833), .S(n22), .Y(n1831) );
  MUX2X1 U1863 ( .B(n1835), .A(n1836), .S(n2259), .Y(n1834) );
  MUX2X1 U1864 ( .B(n1838), .A(n1839), .S(n2259), .Y(n1837) );
  MUX2X1 U1865 ( .B(n1841), .A(n1842), .S(n2259), .Y(n1840) );
  MUX2X1 U1866 ( .B(n1844), .A(n1845), .S(n2259), .Y(n1843) );
  MUX2X1 U1867 ( .B(n1847), .A(n1848), .S(n22), .Y(n1846) );
  MUX2X1 U1868 ( .B(n1850), .A(n1851), .S(n2259), .Y(n1849) );
  MUX2X1 U1869 ( .B(n1853), .A(n1854), .S(n2259), .Y(n1852) );
  MUX2X1 U1870 ( .B(n1856), .A(n1857), .S(n2259), .Y(n1855) );
  MUX2X1 U1871 ( .B(n1859), .A(n1860), .S(n2259), .Y(n1858) );
  MUX2X1 U1872 ( .B(n1862), .A(n1863), .S(n22), .Y(n1861) );
  MUX2X1 U1873 ( .B(n1865), .A(n1866), .S(n20), .Y(n1864) );
  MUX2X1 U1874 ( .B(n1868), .A(n1869), .S(n20), .Y(n1867) );
  MUX2X1 U1875 ( .B(n1871), .A(n1872), .S(n20), .Y(n1870) );
  MUX2X1 U1876 ( .B(n1874), .A(n1875), .S(n20), .Y(n1873) );
  MUX2X1 U1877 ( .B(n1877), .A(n1878), .S(n22), .Y(n1876) );
  MUX2X1 U1878 ( .B(n1880), .A(n1881), .S(n20), .Y(n1879) );
  MUX2X1 U1879 ( .B(n1883), .A(n1884), .S(n20), .Y(n1882) );
  MUX2X1 U1880 ( .B(n1886), .A(n1887), .S(n20), .Y(n1885) );
  MUX2X1 U1881 ( .B(n1889), .A(n1890), .S(n20), .Y(n1888) );
  MUX2X1 U1882 ( .B(n1892), .A(n1893), .S(n22), .Y(n1891) );
  MUX2X1 U1883 ( .B(n1895), .A(n1896), .S(n20), .Y(n1894) );
  MUX2X1 U1884 ( .B(n1898), .A(n1899), .S(n20), .Y(n1897) );
  MUX2X1 U1885 ( .B(n1901), .A(n1902), .S(n20), .Y(n1900) );
  MUX2X1 U1886 ( .B(n1904), .A(n1905), .S(n20), .Y(n1903) );
  MUX2X1 U1887 ( .B(n1907), .A(n1908), .S(n22), .Y(n1906) );
  MUX2X1 U1888 ( .B(n1910), .A(n1911), .S(n20), .Y(n1909) );
  MUX2X1 U1889 ( .B(n1913), .A(n1914), .S(n20), .Y(n1912) );
  MUX2X1 U1890 ( .B(n1916), .A(n1917), .S(n20), .Y(n1915) );
  MUX2X1 U1891 ( .B(n1919), .A(n1920), .S(n20), .Y(n1918) );
  MUX2X1 U1892 ( .B(n1922), .A(n1923), .S(n22), .Y(n1921) );
  MUX2X1 U1893 ( .B(n1925), .A(n1926), .S(n20), .Y(n1924) );
  MUX2X1 U1894 ( .B(n1928), .A(n1929), .S(n20), .Y(n1927) );
  MUX2X1 U1895 ( .B(n1931), .A(n1932), .S(n20), .Y(n1930) );
  MUX2X1 U1896 ( .B(n1934), .A(n1935), .S(n20), .Y(n1933) );
  MUX2X1 U1897 ( .B(n1937), .A(n1938), .S(n22), .Y(n1936) );
  MUX2X1 U1898 ( .B(n1940), .A(n1941), .S(n20), .Y(n1939) );
  MUX2X1 U1899 ( .B(n1943), .A(n1944), .S(n20), .Y(n1942) );
  MUX2X1 U1900 ( .B(n1946), .A(n1947), .S(n20), .Y(n1945) );
  MUX2X1 U1901 ( .B(n1949), .A(n1950), .S(n20), .Y(n1948) );
  MUX2X1 U1902 ( .B(n1952), .A(n1953), .S(n22), .Y(n1951) );
  MUX2X1 U1903 ( .B(n1955), .A(n1956), .S(n20), .Y(n1954) );
  MUX2X1 U1904 ( .B(n1958), .A(n1959), .S(n20), .Y(n1957) );
  MUX2X1 U1905 ( .B(n1961), .A(n1962), .S(n20), .Y(n1960) );
  MUX2X1 U1906 ( .B(n1964), .A(n1965), .S(n20), .Y(n1963) );
  MUX2X1 U1907 ( .B(n1967), .A(n1968), .S(n22), .Y(n1966) );
  MUX2X1 U1908 ( .B(n1970), .A(n1971), .S(n20), .Y(n1969) );
  MUX2X1 U1909 ( .B(n1973), .A(n1974), .S(n20), .Y(n1972) );
  MUX2X1 U1910 ( .B(n1976), .A(n1977), .S(n20), .Y(n1975) );
  MUX2X1 U1911 ( .B(n1979), .A(n1980), .S(n20), .Y(n1978) );
  MUX2X1 U1912 ( .B(n1982), .A(n1983), .S(n22), .Y(n1981) );
  MUX2X1 U1913 ( .B(n1985), .A(n1986), .S(n20), .Y(n1984) );
  MUX2X1 U1914 ( .B(n1988), .A(n1989), .S(n20), .Y(n1987) );
  MUX2X1 U1915 ( .B(n1991), .A(n1992), .S(n20), .Y(n1990) );
  MUX2X1 U1916 ( .B(n1994), .A(n1995), .S(n20), .Y(n1993) );
  MUX2X1 U1917 ( .B(n1997), .A(n1998), .S(n22), .Y(n1996) );
  MUX2X1 U1918 ( .B(n2000), .A(n2001), .S(n20), .Y(n1999) );
  MUX2X1 U1919 ( .B(n2003), .A(n2004), .S(n20), .Y(n2002) );
  MUX2X1 U1920 ( .B(n2006), .A(n2007), .S(n20), .Y(n2005) );
  MUX2X1 U1921 ( .B(n2009), .A(n2010), .S(n20), .Y(n2008) );
  MUX2X1 U1922 ( .B(n2012), .A(n2013), .S(n22), .Y(n2011) );
  MUX2X1 U1923 ( .B(n2015), .A(n2016), .S(n20), .Y(n2014) );
  MUX2X1 U1924 ( .B(n2018), .A(n2019), .S(n20), .Y(n2017) );
  MUX2X1 U1925 ( .B(n2021), .A(n2022), .S(n20), .Y(n2020) );
  MUX2X1 U1926 ( .B(n2024), .A(n2025), .S(n20), .Y(n2023) );
  MUX2X1 U1927 ( .B(n2027), .A(n2028), .S(n22), .Y(n2026) );
  MUX2X1 U1928 ( .B(n2030), .A(n2031), .S(n20), .Y(n2029) );
  MUX2X1 U1929 ( .B(n2033), .A(n2034), .S(n20), .Y(n2032) );
  MUX2X1 U1930 ( .B(n2036), .A(n2037), .S(n20), .Y(n2035) );
  MUX2X1 U1931 ( .B(n2039), .A(n2040), .S(n20), .Y(n2038) );
  MUX2X1 U1932 ( .B(n2042), .A(n2043), .S(n22), .Y(n2041) );
  MUX2X1 U1933 ( .B(n2045), .A(n2046), .S(n20), .Y(n2044) );
  MUX2X1 U1934 ( .B(n2048), .A(n2049), .S(n20), .Y(n2047) );
  MUX2X1 U1935 ( .B(n2051), .A(n2052), .S(n20), .Y(n2050) );
  MUX2X1 U1936 ( .B(n2054), .A(n2055), .S(n20), .Y(n2053) );
  MUX2X1 U1937 ( .B(n2057), .A(n2058), .S(n22), .Y(n2056) );
  MUX2X1 U1938 ( .B(n2060), .A(n2061), .S(n20), .Y(n2059) );
  MUX2X1 U1939 ( .B(n2063), .A(n2064), .S(n20), .Y(n2062) );
  MUX2X1 U1940 ( .B(n2066), .A(n2067), .S(n20), .Y(n2065) );
  MUX2X1 U1941 ( .B(n2069), .A(n2070), .S(n20), .Y(n2068) );
  MUX2X1 U1942 ( .B(n2072), .A(n2073), .S(n22), .Y(n2071) );
  MUX2X1 U1943 ( .B(n2075), .A(n2076), .S(n20), .Y(n2074) );
  MUX2X1 U1944 ( .B(n2078), .A(n2079), .S(n20), .Y(n2077) );
  MUX2X1 U1945 ( .B(n2081), .A(n2082), .S(n20), .Y(n2080) );
  MUX2X1 U1946 ( .B(n2084), .A(n2085), .S(n20), .Y(n2083) );
  MUX2X1 U1947 ( .B(n2087), .A(n2088), .S(n22), .Y(n2086) );
  MUX2X1 U1948 ( .B(n2090), .A(n2091), .S(n20), .Y(n2089) );
  MUX2X1 U1949 ( .B(n2093), .A(n2094), .S(n20), .Y(n2092) );
  MUX2X1 U1950 ( .B(n2096), .A(n2097), .S(n20), .Y(n2095) );
  MUX2X1 U1951 ( .B(n2099), .A(n2100), .S(n20), .Y(n2098) );
  MUX2X1 U1952 ( .B(n2102), .A(n2103), .S(n22), .Y(n2101) );
  MUX2X1 U1953 ( .B(n2105), .A(n2106), .S(n20), .Y(n2104) );
  MUX2X1 U1954 ( .B(n2108), .A(n2109), .S(n20), .Y(n2107) );
  MUX2X1 U1955 ( .B(n2111), .A(n2112), .S(n20), .Y(n2110) );
  MUX2X1 U1956 ( .B(n2114), .A(n2115), .S(n20), .Y(n2113) );
  MUX2X1 U1957 ( .B(n2117), .A(n2118), .S(n22), .Y(n2116) );
  MUX2X1 U1958 ( .B(n2120), .A(n2121), .S(n20), .Y(n2119) );
  MUX2X1 U1959 ( .B(n2123), .A(n2124), .S(n20), .Y(n2122) );
  MUX2X1 U1960 ( .B(n2126), .A(n2127), .S(n20), .Y(n2125) );
  MUX2X1 U1961 ( .B(n2129), .A(n2130), .S(n20), .Y(n2128) );
  MUX2X1 U1962 ( .B(n2132), .A(n2133), .S(n22), .Y(n2131) );
  MUX2X1 U1963 ( .B(n2135), .A(n2136), .S(n20), .Y(n2134) );
  MUX2X1 U1964 ( .B(n2138), .A(n2139), .S(n20), .Y(n2137) );
  MUX2X1 U1965 ( .B(n2141), .A(n2142), .S(n20), .Y(n2140) );
  MUX2X1 U1966 ( .B(n2144), .A(n2145), .S(n20), .Y(n2143) );
  MUX2X1 U1967 ( .B(n2147), .A(n2148), .S(n22), .Y(n2146) );
  MUX2X1 U1968 ( .B(n2150), .A(n2151), .S(n20), .Y(n2149) );
  MUX2X1 U1969 ( .B(n2153), .A(n2154), .S(n20), .Y(n2152) );
  MUX2X1 U1970 ( .B(n2156), .A(n2157), .S(n20), .Y(n2155) );
  MUX2X1 U1971 ( .B(n2159), .A(n2160), .S(n20), .Y(n2158) );
  MUX2X1 U1972 ( .B(n2162), .A(n2163), .S(n22), .Y(n2161) );
  MUX2X1 U1973 ( .B(n2165), .A(n2166), .S(n20), .Y(n2164) );
  MUX2X1 U1974 ( .B(n2168), .A(n2169), .S(n20), .Y(n2167) );
  MUX2X1 U1975 ( .B(n2171), .A(n2172), .S(n20), .Y(n2170) );
  MUX2X1 U1976 ( .B(n2174), .A(n2175), .S(n20), .Y(n2173) );
  MUX2X1 U1977 ( .B(n2177), .A(n2178), .S(n22), .Y(n2176) );
  MUX2X1 U1978 ( .B(n2180), .A(n2181), .S(n20), .Y(n2179) );
  MUX2X1 U1979 ( .B(n2183), .A(n2184), .S(n2259), .Y(n2182) );
  MUX2X1 U1980 ( .B(n2186), .A(n2187), .S(n2258), .Y(n2185) );
  MUX2X1 U1981 ( .B(n2189), .A(n2190), .S(n20), .Y(n2188) );
  MUX2X1 U1982 ( .B(n2192), .A(n2193), .S(n22), .Y(n2191) );
  MUX2X1 U1983 ( .B(n2195), .A(n2196), .S(n20), .Y(n2194) );
  MUX2X1 U1984 ( .B(n2198), .A(n2199), .S(n20), .Y(n2197) );
  MUX2X1 U1985 ( .B(n2201), .A(n2202), .S(n20), .Y(n2200) );
  MUX2X1 U1986 ( .B(n2204), .A(n2205), .S(n20), .Y(n2203) );
  MUX2X1 U1987 ( .B(n2207), .A(n2208), .S(n22), .Y(n2206) );
  MUX2X1 U1988 ( .B(n2210), .A(n2211), .S(n20), .Y(n2209) );
  MUX2X1 U1989 ( .B(n2213), .A(n2214), .S(n20), .Y(n2212) );
  MUX2X1 U1990 ( .B(n2216), .A(n2217), .S(n2259), .Y(n2215) );
  MUX2X1 U1991 ( .B(n2219), .A(n2220), .S(n2258), .Y(n2218) );
  MUX2X1 U1992 ( .B(n2222), .A(n2223), .S(n22), .Y(n2221) );
  MUX2X1 U1993 ( .B(fifo_array[480]), .A(fifo_array[496]), .S(n19), .Y(n1746)
         );
  MUX2X1 U1994 ( .B(fifo_array[448]), .A(fifo_array[464]), .S(n19), .Y(n1745)
         );
  MUX2X1 U1995 ( .B(fifo_array[416]), .A(fifo_array[432]), .S(n2311), .Y(n1749) );
  MUX2X1 U1996 ( .B(fifo_array[384]), .A(fifo_array[400]), .S(n2257), .Y(n1748) );
  MUX2X1 U1997 ( .B(n1747), .A(n1744), .S(n21), .Y(n1758) );
  MUX2X1 U1998 ( .B(fifo_array[352]), .A(fifo_array[368]), .S(n2241), .Y(n1752) );
  MUX2X1 U1999 ( .B(fifo_array[320]), .A(fifo_array[336]), .S(n2241), .Y(n1751) );
  MUX2X1 U2000 ( .B(fifo_array[288]), .A(fifo_array[304]), .S(n2241), .Y(n1755) );
  MUX2X1 U2001 ( .B(fifo_array[256]), .A(fifo_array[272]), .S(n2241), .Y(n1754) );
  MUX2X1 U2002 ( .B(n1753), .A(n1750), .S(n21), .Y(n1757) );
  MUX2X1 U2003 ( .B(fifo_array[224]), .A(fifo_array[240]), .S(n2241), .Y(n1761) );
  MUX2X1 U2004 ( .B(fifo_array[192]), .A(fifo_array[208]), .S(n2241), .Y(n1760) );
  MUX2X1 U2005 ( .B(fifo_array[160]), .A(fifo_array[176]), .S(n2241), .Y(n1764) );
  MUX2X1 U2006 ( .B(fifo_array[128]), .A(fifo_array[144]), .S(n2241), .Y(n1763) );
  MUX2X1 U2007 ( .B(n1762), .A(n1759), .S(n21), .Y(n1773) );
  MUX2X1 U2008 ( .B(fifo_array[96]), .A(fifo_array[112]), .S(n2241), .Y(n1767)
         );
  MUX2X1 U2009 ( .B(fifo_array[64]), .A(fifo_array[80]), .S(n2241), .Y(n1766)
         );
  MUX2X1 U2010 ( .B(fifo_array[32]), .A(fifo_array[48]), .S(n2241), .Y(n1770)
         );
  MUX2X1 U2011 ( .B(fifo_array[0]), .A(fifo_array[16]), .S(n2241), .Y(n1769)
         );
  MUX2X1 U2012 ( .B(n1768), .A(n1765), .S(n21), .Y(n1772) );
  MUX2X1 U2013 ( .B(n1771), .A(n1756), .S(n23), .Y(n2224) );
  MUX2X1 U2014 ( .B(fifo_array[481]), .A(fifo_array[497]), .S(n2242), .Y(n1776) );
  MUX2X1 U2015 ( .B(fifo_array[449]), .A(fifo_array[465]), .S(n2242), .Y(n1775) );
  MUX2X1 U2016 ( .B(fifo_array[417]), .A(fifo_array[433]), .S(n2242), .Y(n1779) );
  MUX2X1 U2017 ( .B(fifo_array[385]), .A(fifo_array[401]), .S(n2242), .Y(n1778) );
  MUX2X1 U2018 ( .B(n1777), .A(n1774), .S(n21), .Y(n1788) );
  MUX2X1 U2019 ( .B(fifo_array[353]), .A(fifo_array[369]), .S(n2242), .Y(n1782) );
  MUX2X1 U2020 ( .B(fifo_array[321]), .A(fifo_array[337]), .S(n2242), .Y(n1781) );
  MUX2X1 U2021 ( .B(fifo_array[289]), .A(fifo_array[305]), .S(n2242), .Y(n1785) );
  MUX2X1 U2022 ( .B(fifo_array[257]), .A(fifo_array[273]), .S(n2242), .Y(n1784) );
  MUX2X1 U2023 ( .B(n1783), .A(n1780), .S(n21), .Y(n1787) );
  MUX2X1 U2024 ( .B(fifo_array[225]), .A(fifo_array[241]), .S(n2242), .Y(n1791) );
  MUX2X1 U2025 ( .B(fifo_array[193]), .A(fifo_array[209]), .S(n2242), .Y(n1790) );
  MUX2X1 U2026 ( .B(fifo_array[161]), .A(fifo_array[177]), .S(n2242), .Y(n1794) );
  MUX2X1 U2027 ( .B(fifo_array[129]), .A(fifo_array[145]), .S(n2242), .Y(n1793) );
  MUX2X1 U2028 ( .B(n1792), .A(n1789), .S(n21), .Y(n1803) );
  MUX2X1 U2029 ( .B(fifo_array[97]), .A(fifo_array[113]), .S(n2243), .Y(n1797)
         );
  MUX2X1 U2030 ( .B(fifo_array[65]), .A(fifo_array[81]), .S(n2243), .Y(n1796)
         );
  MUX2X1 U2031 ( .B(fifo_array[33]), .A(fifo_array[49]), .S(n2243), .Y(n1800)
         );
  MUX2X1 U2032 ( .B(fifo_array[1]), .A(fifo_array[17]), .S(n2243), .Y(n1799)
         );
  MUX2X1 U2033 ( .B(n1798), .A(n1795), .S(n21), .Y(n1802) );
  MUX2X1 U2034 ( .B(n1801), .A(n1786), .S(n23), .Y(n2225) );
  MUX2X1 U2035 ( .B(fifo_array[482]), .A(fifo_array[498]), .S(n2243), .Y(n1806) );
  MUX2X1 U2036 ( .B(fifo_array[450]), .A(fifo_array[466]), .S(n2243), .Y(n1805) );
  MUX2X1 U2037 ( .B(fifo_array[418]), .A(fifo_array[434]), .S(n2243), .Y(n1809) );
  MUX2X1 U2038 ( .B(fifo_array[386]), .A(fifo_array[402]), .S(n2243), .Y(n1808) );
  MUX2X1 U2039 ( .B(n1807), .A(n1804), .S(n21), .Y(n1818) );
  MUX2X1 U2040 ( .B(fifo_array[354]), .A(fifo_array[370]), .S(n2243), .Y(n1812) );
  MUX2X1 U2041 ( .B(fifo_array[322]), .A(fifo_array[338]), .S(n2243), .Y(n1811) );
  MUX2X1 U2042 ( .B(fifo_array[290]), .A(fifo_array[306]), .S(n2243), .Y(n1815) );
  MUX2X1 U2043 ( .B(fifo_array[258]), .A(fifo_array[274]), .S(n2243), .Y(n1814) );
  MUX2X1 U2044 ( .B(n1813), .A(n1810), .S(n21), .Y(n1817) );
  MUX2X1 U2045 ( .B(fifo_array[226]), .A(fifo_array[242]), .S(n2244), .Y(n1821) );
  MUX2X1 U2046 ( .B(fifo_array[194]), .A(fifo_array[210]), .S(n2244), .Y(n1820) );
  MUX2X1 U2047 ( .B(fifo_array[162]), .A(fifo_array[178]), .S(n2244), .Y(n1824) );
  MUX2X1 U2048 ( .B(fifo_array[130]), .A(fifo_array[146]), .S(n2244), .Y(n1823) );
  MUX2X1 U2049 ( .B(n1822), .A(n1819), .S(n21), .Y(n1833) );
  MUX2X1 U2050 ( .B(fifo_array[98]), .A(fifo_array[114]), .S(n2244), .Y(n1827)
         );
  MUX2X1 U2051 ( .B(fifo_array[66]), .A(fifo_array[82]), .S(n2244), .Y(n1826)
         );
  MUX2X1 U2052 ( .B(fifo_array[34]), .A(fifo_array[50]), .S(n2244), .Y(n1830)
         );
  MUX2X1 U2053 ( .B(fifo_array[2]), .A(fifo_array[18]), .S(n2244), .Y(n1829)
         );
  MUX2X1 U2054 ( .B(n1828), .A(n1825), .S(n21), .Y(n1832) );
  MUX2X1 U2055 ( .B(n1831), .A(n1816), .S(n23), .Y(n2226) );
  MUX2X1 U2056 ( .B(fifo_array[483]), .A(fifo_array[499]), .S(n2244), .Y(n1836) );
  MUX2X1 U2057 ( .B(fifo_array[451]), .A(fifo_array[467]), .S(n2244), .Y(n1835) );
  MUX2X1 U2058 ( .B(fifo_array[419]), .A(fifo_array[435]), .S(n2244), .Y(n1839) );
  MUX2X1 U2059 ( .B(fifo_array[387]), .A(fifo_array[403]), .S(n2244), .Y(n1838) );
  MUX2X1 U2060 ( .B(n1837), .A(n1834), .S(n21), .Y(n1848) );
  MUX2X1 U2061 ( .B(fifo_array[355]), .A(fifo_array[371]), .S(n2245), .Y(n1842) );
  MUX2X1 U2062 ( .B(fifo_array[323]), .A(fifo_array[339]), .S(n2245), .Y(n1841) );
  MUX2X1 U2063 ( .B(fifo_array[291]), .A(fifo_array[307]), .S(n2245), .Y(n1845) );
  MUX2X1 U2064 ( .B(fifo_array[259]), .A(fifo_array[275]), .S(n2245), .Y(n1844) );
  MUX2X1 U2065 ( .B(n1843), .A(n1840), .S(n21), .Y(n1847) );
  MUX2X1 U2066 ( .B(fifo_array[227]), .A(fifo_array[243]), .S(n2245), .Y(n1851) );
  MUX2X1 U2067 ( .B(fifo_array[195]), .A(fifo_array[211]), .S(n2245), .Y(n1850) );
  MUX2X1 U2068 ( .B(fifo_array[163]), .A(fifo_array[179]), .S(n2245), .Y(n1854) );
  MUX2X1 U2069 ( .B(fifo_array[131]), .A(fifo_array[147]), .S(n2245), .Y(n1853) );
  MUX2X1 U2070 ( .B(n1852), .A(n1849), .S(n21), .Y(n1863) );
  MUX2X1 U2071 ( .B(fifo_array[99]), .A(fifo_array[115]), .S(n2245), .Y(n1857)
         );
  MUX2X1 U2072 ( .B(fifo_array[67]), .A(fifo_array[83]), .S(n2245), .Y(n1856)
         );
  MUX2X1 U2073 ( .B(fifo_array[35]), .A(fifo_array[51]), .S(n2245), .Y(n1860)
         );
  MUX2X1 U2074 ( .B(fifo_array[3]), .A(fifo_array[19]), .S(n2245), .Y(n1859)
         );
  MUX2X1 U2075 ( .B(n1858), .A(n1855), .S(n21), .Y(n1862) );
  MUX2X1 U2076 ( .B(n1861), .A(n1846), .S(n23), .Y(n2227) );
  MUX2X1 U2077 ( .B(fifo_array[484]), .A(fifo_array[500]), .S(n2246), .Y(n1866) );
  MUX2X1 U2078 ( .B(fifo_array[452]), .A(fifo_array[468]), .S(n2246), .Y(n1865) );
  MUX2X1 U2079 ( .B(fifo_array[420]), .A(fifo_array[436]), .S(n2246), .Y(n1869) );
  MUX2X1 U2080 ( .B(fifo_array[388]), .A(fifo_array[404]), .S(n2246), .Y(n1868) );
  MUX2X1 U2081 ( .B(n1867), .A(n1864), .S(n21), .Y(n1878) );
  MUX2X1 U2082 ( .B(fifo_array[356]), .A(fifo_array[372]), .S(n2246), .Y(n1872) );
  MUX2X1 U2083 ( .B(fifo_array[324]), .A(fifo_array[340]), .S(n2246), .Y(n1871) );
  MUX2X1 U2084 ( .B(fifo_array[292]), .A(fifo_array[308]), .S(n2246), .Y(n1875) );
  MUX2X1 U2085 ( .B(fifo_array[260]), .A(fifo_array[276]), .S(n2246), .Y(n1874) );
  MUX2X1 U2086 ( .B(n1873), .A(n1870), .S(n21), .Y(n1877) );
  MUX2X1 U2087 ( .B(fifo_array[228]), .A(fifo_array[244]), .S(n2246), .Y(n1881) );
  MUX2X1 U2088 ( .B(fifo_array[196]), .A(fifo_array[212]), .S(n2246), .Y(n1880) );
  MUX2X1 U2089 ( .B(fifo_array[164]), .A(fifo_array[180]), .S(n2246), .Y(n1884) );
  MUX2X1 U2090 ( .B(fifo_array[132]), .A(fifo_array[148]), .S(n2246), .Y(n1883) );
  MUX2X1 U2091 ( .B(n1882), .A(n1879), .S(n21), .Y(n1893) );
  MUX2X1 U2092 ( .B(fifo_array[100]), .A(fifo_array[116]), .S(n2247), .Y(n1887) );
  MUX2X1 U2093 ( .B(fifo_array[68]), .A(fifo_array[84]), .S(n2247), .Y(n1886)
         );
  MUX2X1 U2094 ( .B(fifo_array[36]), .A(fifo_array[52]), .S(n2247), .Y(n1890)
         );
  MUX2X1 U2095 ( .B(fifo_array[4]), .A(fifo_array[20]), .S(n2247), .Y(n1889)
         );
  MUX2X1 U2096 ( .B(n1888), .A(n1885), .S(n21), .Y(n1892) );
  MUX2X1 U2097 ( .B(n1891), .A(n1876), .S(n23), .Y(n2228) );
  MUX2X1 U2098 ( .B(fifo_array[485]), .A(fifo_array[501]), .S(n2247), .Y(n1896) );
  MUX2X1 U2099 ( .B(fifo_array[453]), .A(fifo_array[469]), .S(n2247), .Y(n1895) );
  MUX2X1 U2100 ( .B(fifo_array[421]), .A(fifo_array[437]), .S(n2247), .Y(n1899) );
  MUX2X1 U2101 ( .B(fifo_array[389]), .A(fifo_array[405]), .S(n2247), .Y(n1898) );
  MUX2X1 U2102 ( .B(n1897), .A(n1894), .S(n21), .Y(n1908) );
  MUX2X1 U2103 ( .B(fifo_array[357]), .A(fifo_array[373]), .S(n2247), .Y(n1902) );
  MUX2X1 U2104 ( .B(fifo_array[325]), .A(fifo_array[341]), .S(n2247), .Y(n1901) );
  MUX2X1 U2105 ( .B(fifo_array[293]), .A(fifo_array[309]), .S(n2247), .Y(n1905) );
  MUX2X1 U2106 ( .B(fifo_array[261]), .A(fifo_array[277]), .S(n2247), .Y(n1904) );
  MUX2X1 U2107 ( .B(n1903), .A(n1900), .S(n21), .Y(n1907) );
  MUX2X1 U2108 ( .B(fifo_array[229]), .A(fifo_array[245]), .S(n2248), .Y(n1911) );
  MUX2X1 U2109 ( .B(fifo_array[197]), .A(fifo_array[213]), .S(n2248), .Y(n1910) );
  MUX2X1 U2110 ( .B(fifo_array[165]), .A(fifo_array[181]), .S(n2248), .Y(n1914) );
  MUX2X1 U2111 ( .B(fifo_array[133]), .A(fifo_array[149]), .S(n2248), .Y(n1913) );
  MUX2X1 U2112 ( .B(n1912), .A(n1909), .S(n21), .Y(n1923) );
  MUX2X1 U2113 ( .B(fifo_array[101]), .A(fifo_array[117]), .S(n2248), .Y(n1917) );
  MUX2X1 U2114 ( .B(fifo_array[69]), .A(fifo_array[85]), .S(n2248), .Y(n1916)
         );
  MUX2X1 U2115 ( .B(fifo_array[37]), .A(fifo_array[53]), .S(n2248), .Y(n1920)
         );
  MUX2X1 U2116 ( .B(fifo_array[5]), .A(fifo_array[21]), .S(n2248), .Y(n1919)
         );
  MUX2X1 U2117 ( .B(n1918), .A(n1915), .S(n21), .Y(n1922) );
  MUX2X1 U2118 ( .B(n1921), .A(n1906), .S(n23), .Y(n2229) );
  MUX2X1 U2119 ( .B(fifo_array[486]), .A(fifo_array[502]), .S(n2248), .Y(n1926) );
  MUX2X1 U2120 ( .B(fifo_array[454]), .A(fifo_array[470]), .S(n2248), .Y(n1925) );
  MUX2X1 U2121 ( .B(fifo_array[422]), .A(fifo_array[438]), .S(n2248), .Y(n1929) );
  MUX2X1 U2122 ( .B(fifo_array[390]), .A(fifo_array[406]), .S(n2248), .Y(n1928) );
  MUX2X1 U2123 ( .B(n1927), .A(n1924), .S(n21), .Y(n1938) );
  MUX2X1 U2124 ( .B(fifo_array[358]), .A(fifo_array[374]), .S(n2249), .Y(n1932) );
  MUX2X1 U2125 ( .B(fifo_array[326]), .A(fifo_array[342]), .S(n2249), .Y(n1931) );
  MUX2X1 U2126 ( .B(fifo_array[294]), .A(fifo_array[310]), .S(n2249), .Y(n1935) );
  MUX2X1 U2127 ( .B(fifo_array[262]), .A(fifo_array[278]), .S(n2249), .Y(n1934) );
  MUX2X1 U2128 ( .B(n1933), .A(n1930), .S(n21), .Y(n1937) );
  MUX2X1 U2129 ( .B(fifo_array[230]), .A(fifo_array[246]), .S(n2249), .Y(n1941) );
  MUX2X1 U2130 ( .B(fifo_array[198]), .A(fifo_array[214]), .S(n2249), .Y(n1940) );
  MUX2X1 U2131 ( .B(fifo_array[166]), .A(fifo_array[182]), .S(n2249), .Y(n1944) );
  MUX2X1 U2132 ( .B(fifo_array[134]), .A(fifo_array[150]), .S(n2249), .Y(n1943) );
  MUX2X1 U2133 ( .B(n1942), .A(n1939), .S(n21), .Y(n1953) );
  MUX2X1 U2134 ( .B(fifo_array[102]), .A(fifo_array[118]), .S(n2249), .Y(n1947) );
  MUX2X1 U2135 ( .B(fifo_array[70]), .A(fifo_array[86]), .S(n2249), .Y(n1946)
         );
  MUX2X1 U2136 ( .B(fifo_array[38]), .A(fifo_array[54]), .S(n2249), .Y(n1950)
         );
  MUX2X1 U2137 ( .B(fifo_array[6]), .A(fifo_array[22]), .S(n2249), .Y(n1949)
         );
  MUX2X1 U2138 ( .B(n1948), .A(n1945), .S(n21), .Y(n1952) );
  MUX2X1 U2139 ( .B(n1951), .A(n1936), .S(n23), .Y(n2230) );
  MUX2X1 U2140 ( .B(fifo_array[487]), .A(fifo_array[503]), .S(n2250), .Y(n1956) );
  MUX2X1 U2141 ( .B(fifo_array[455]), .A(fifo_array[471]), .S(n2250), .Y(n1955) );
  MUX2X1 U2142 ( .B(fifo_array[423]), .A(fifo_array[439]), .S(n2250), .Y(n1959) );
  MUX2X1 U2143 ( .B(fifo_array[391]), .A(fifo_array[407]), .S(n2250), .Y(n1958) );
  MUX2X1 U2144 ( .B(n1957), .A(n1954), .S(n21), .Y(n1968) );
  MUX2X1 U2145 ( .B(fifo_array[359]), .A(fifo_array[375]), .S(n2250), .Y(n1962) );
  MUX2X1 U2146 ( .B(fifo_array[327]), .A(fifo_array[343]), .S(n2250), .Y(n1961) );
  MUX2X1 U2147 ( .B(fifo_array[295]), .A(fifo_array[311]), .S(n2250), .Y(n1965) );
  MUX2X1 U2148 ( .B(fifo_array[263]), .A(fifo_array[279]), .S(n2250), .Y(n1964) );
  MUX2X1 U2149 ( .B(n1963), .A(n1960), .S(n21), .Y(n1967) );
  MUX2X1 U2150 ( .B(fifo_array[231]), .A(fifo_array[247]), .S(n2250), .Y(n1971) );
  MUX2X1 U2151 ( .B(fifo_array[199]), .A(fifo_array[215]), .S(n2250), .Y(n1970) );
  MUX2X1 U2152 ( .B(fifo_array[167]), .A(fifo_array[183]), .S(n2250), .Y(n1974) );
  MUX2X1 U2153 ( .B(fifo_array[135]), .A(fifo_array[151]), .S(n2250), .Y(n1973) );
  MUX2X1 U2154 ( .B(n1972), .A(n1969), .S(n21), .Y(n1983) );
  MUX2X1 U2155 ( .B(fifo_array[103]), .A(fifo_array[119]), .S(n2251), .Y(n1977) );
  MUX2X1 U2156 ( .B(fifo_array[71]), .A(fifo_array[87]), .S(n2251), .Y(n1976)
         );
  MUX2X1 U2157 ( .B(fifo_array[39]), .A(fifo_array[55]), .S(n2251), .Y(n1980)
         );
  MUX2X1 U2158 ( .B(fifo_array[7]), .A(fifo_array[23]), .S(n2251), .Y(n1979)
         );
  MUX2X1 U2159 ( .B(n1978), .A(n1975), .S(n21), .Y(n1982) );
  MUX2X1 U2160 ( .B(n1981), .A(n1966), .S(n23), .Y(n2231) );
  MUX2X1 U2161 ( .B(fifo_array[488]), .A(fifo_array[504]), .S(n2251), .Y(n1986) );
  MUX2X1 U2162 ( .B(fifo_array[456]), .A(fifo_array[472]), .S(n2251), .Y(n1985) );
  MUX2X1 U2163 ( .B(fifo_array[424]), .A(fifo_array[440]), .S(n2251), .Y(n1989) );
  MUX2X1 U2164 ( .B(fifo_array[392]), .A(fifo_array[408]), .S(n2251), .Y(n1988) );
  MUX2X1 U2165 ( .B(n1987), .A(n1984), .S(n21), .Y(n1998) );
  MUX2X1 U2166 ( .B(fifo_array[360]), .A(fifo_array[376]), .S(n2251), .Y(n1992) );
  MUX2X1 U2167 ( .B(fifo_array[328]), .A(fifo_array[344]), .S(n2251), .Y(n1991) );
  MUX2X1 U2168 ( .B(fifo_array[296]), .A(fifo_array[312]), .S(n2251), .Y(n1995) );
  MUX2X1 U2169 ( .B(fifo_array[264]), .A(fifo_array[280]), .S(n2251), .Y(n1994) );
  MUX2X1 U2170 ( .B(n1993), .A(n1990), .S(n21), .Y(n1997) );
  MUX2X1 U2171 ( .B(fifo_array[232]), .A(fifo_array[248]), .S(n2252), .Y(n2001) );
  MUX2X1 U2172 ( .B(fifo_array[200]), .A(fifo_array[216]), .S(n2252), .Y(n2000) );
  MUX2X1 U2173 ( .B(fifo_array[168]), .A(fifo_array[184]), .S(n2252), .Y(n2004) );
  MUX2X1 U2174 ( .B(fifo_array[136]), .A(fifo_array[152]), .S(n2252), .Y(n2003) );
  MUX2X1 U2175 ( .B(n2002), .A(n1999), .S(n21), .Y(n2013) );
  MUX2X1 U2176 ( .B(fifo_array[104]), .A(fifo_array[120]), .S(n2252), .Y(n2007) );
  MUX2X1 U2177 ( .B(fifo_array[72]), .A(fifo_array[88]), .S(n2252), .Y(n2006)
         );
  MUX2X1 U2178 ( .B(fifo_array[40]), .A(fifo_array[56]), .S(n2252), .Y(n2010)
         );
  MUX2X1 U2179 ( .B(fifo_array[8]), .A(fifo_array[24]), .S(n2252), .Y(n2009)
         );
  MUX2X1 U2180 ( .B(n2008), .A(n2005), .S(n21), .Y(n2012) );
  MUX2X1 U2181 ( .B(n2011), .A(n1996), .S(n23), .Y(n2232) );
  MUX2X1 U2182 ( .B(fifo_array[489]), .A(fifo_array[505]), .S(n2252), .Y(n2016) );
  MUX2X1 U2183 ( .B(fifo_array[457]), .A(fifo_array[473]), .S(n2252), .Y(n2015) );
  MUX2X1 U2184 ( .B(fifo_array[425]), .A(fifo_array[441]), .S(n2252), .Y(n2019) );
  MUX2X1 U2185 ( .B(fifo_array[393]), .A(fifo_array[409]), .S(n2252), .Y(n2018) );
  MUX2X1 U2186 ( .B(n2017), .A(n2014), .S(n21), .Y(n2028) );
  MUX2X1 U2187 ( .B(fifo_array[361]), .A(fifo_array[377]), .S(n2253), .Y(n2022) );
  MUX2X1 U2188 ( .B(fifo_array[329]), .A(fifo_array[345]), .S(n2253), .Y(n2021) );
  MUX2X1 U2189 ( .B(fifo_array[297]), .A(fifo_array[313]), .S(n2253), .Y(n2025) );
  MUX2X1 U2190 ( .B(fifo_array[265]), .A(fifo_array[281]), .S(n2253), .Y(n2024) );
  MUX2X1 U2191 ( .B(n2023), .A(n2020), .S(n21), .Y(n2027) );
  MUX2X1 U2192 ( .B(fifo_array[233]), .A(fifo_array[249]), .S(n2253), .Y(n2031) );
  MUX2X1 U2193 ( .B(fifo_array[201]), .A(fifo_array[217]), .S(n2253), .Y(n2030) );
  MUX2X1 U2194 ( .B(fifo_array[169]), .A(fifo_array[185]), .S(n2253), .Y(n2034) );
  MUX2X1 U2195 ( .B(fifo_array[137]), .A(fifo_array[153]), .S(n2253), .Y(n2033) );
  MUX2X1 U2196 ( .B(n2032), .A(n2029), .S(n21), .Y(n2043) );
  MUX2X1 U2197 ( .B(fifo_array[105]), .A(fifo_array[121]), .S(n2253), .Y(n2037) );
  MUX2X1 U2198 ( .B(fifo_array[73]), .A(fifo_array[89]), .S(n2253), .Y(n2036)
         );
  MUX2X1 U2199 ( .B(fifo_array[41]), .A(fifo_array[57]), .S(n2253), .Y(n2040)
         );
  MUX2X1 U2200 ( .B(fifo_array[9]), .A(fifo_array[25]), .S(n2253), .Y(n2039)
         );
  MUX2X1 U2201 ( .B(n2038), .A(n2035), .S(n21), .Y(n2042) );
  MUX2X1 U2202 ( .B(n2041), .A(n2026), .S(n23), .Y(n2233) );
  MUX2X1 U2203 ( .B(fifo_array[490]), .A(fifo_array[506]), .S(n2254), .Y(n2046) );
  MUX2X1 U2204 ( .B(fifo_array[458]), .A(fifo_array[474]), .S(n2254), .Y(n2045) );
  MUX2X1 U2205 ( .B(fifo_array[426]), .A(fifo_array[442]), .S(n2254), .Y(n2049) );
  MUX2X1 U2206 ( .B(fifo_array[394]), .A(fifo_array[410]), .S(n2254), .Y(n2048) );
  MUX2X1 U2207 ( .B(n2047), .A(n2044), .S(n21), .Y(n2058) );
  MUX2X1 U2208 ( .B(fifo_array[362]), .A(fifo_array[378]), .S(n2254), .Y(n2052) );
  MUX2X1 U2209 ( .B(fifo_array[330]), .A(fifo_array[346]), .S(n2254), .Y(n2051) );
  MUX2X1 U2210 ( .B(fifo_array[298]), .A(fifo_array[314]), .S(n2254), .Y(n2055) );
  MUX2X1 U2211 ( .B(fifo_array[266]), .A(fifo_array[282]), .S(n2254), .Y(n2054) );
  MUX2X1 U2212 ( .B(n2053), .A(n2050), .S(n21), .Y(n2057) );
  MUX2X1 U2213 ( .B(fifo_array[234]), .A(fifo_array[250]), .S(n2254), .Y(n2061) );
  MUX2X1 U2214 ( .B(fifo_array[202]), .A(fifo_array[218]), .S(n2254), .Y(n2060) );
  MUX2X1 U2215 ( .B(fifo_array[170]), .A(fifo_array[186]), .S(n2254), .Y(n2064) );
  MUX2X1 U2216 ( .B(fifo_array[138]), .A(fifo_array[154]), .S(n2254), .Y(n2063) );
  MUX2X1 U2217 ( .B(n2062), .A(n2059), .S(n21), .Y(n2073) );
  MUX2X1 U2218 ( .B(fifo_array[106]), .A(fifo_array[122]), .S(n2255), .Y(n2067) );
  MUX2X1 U2219 ( .B(fifo_array[74]), .A(fifo_array[90]), .S(n2255), .Y(n2066)
         );
  MUX2X1 U2220 ( .B(fifo_array[42]), .A(fifo_array[58]), .S(n2255), .Y(n2070)
         );
  MUX2X1 U2221 ( .B(fifo_array[10]), .A(fifo_array[26]), .S(n2255), .Y(n2069)
         );
  MUX2X1 U2222 ( .B(n2068), .A(n2065), .S(n21), .Y(n2072) );
  MUX2X1 U2223 ( .B(n2071), .A(n2056), .S(n23), .Y(n2234) );
  MUX2X1 U2224 ( .B(fifo_array[491]), .A(fifo_array[507]), .S(n2255), .Y(n2076) );
  MUX2X1 U2225 ( .B(fifo_array[459]), .A(fifo_array[475]), .S(n2255), .Y(n2075) );
  MUX2X1 U2226 ( .B(fifo_array[427]), .A(fifo_array[443]), .S(n2255), .Y(n2079) );
  MUX2X1 U2227 ( .B(fifo_array[395]), .A(fifo_array[411]), .S(n2255), .Y(n2078) );
  MUX2X1 U2228 ( .B(n2077), .A(n2074), .S(n21), .Y(n2088) );
  MUX2X1 U2229 ( .B(fifo_array[363]), .A(fifo_array[379]), .S(n2255), .Y(n2082) );
  MUX2X1 U2230 ( .B(fifo_array[331]), .A(fifo_array[347]), .S(n2255), .Y(n2081) );
  MUX2X1 U2231 ( .B(fifo_array[299]), .A(fifo_array[315]), .S(n2255), .Y(n2085) );
  MUX2X1 U2232 ( .B(fifo_array[267]), .A(fifo_array[283]), .S(n2255), .Y(n2084) );
  MUX2X1 U2233 ( .B(n2083), .A(n2080), .S(n21), .Y(n2087) );
  MUX2X1 U2234 ( .B(fifo_array[235]), .A(fifo_array[251]), .S(n2256), .Y(n2091) );
  MUX2X1 U2235 ( .B(fifo_array[203]), .A(fifo_array[219]), .S(n2256), .Y(n2090) );
  MUX2X1 U2236 ( .B(fifo_array[171]), .A(fifo_array[187]), .S(n2256), .Y(n2094) );
  MUX2X1 U2237 ( .B(fifo_array[139]), .A(fifo_array[155]), .S(n2256), .Y(n2093) );
  MUX2X1 U2238 ( .B(n2092), .A(n2089), .S(n21), .Y(n2103) );
  MUX2X1 U2239 ( .B(fifo_array[107]), .A(fifo_array[123]), .S(n2256), .Y(n2097) );
  MUX2X1 U2240 ( .B(fifo_array[75]), .A(fifo_array[91]), .S(n2256), .Y(n2096)
         );
  MUX2X1 U2241 ( .B(fifo_array[43]), .A(fifo_array[59]), .S(n2256), .Y(n2100)
         );
  MUX2X1 U2242 ( .B(fifo_array[11]), .A(fifo_array[27]), .S(n2256), .Y(n2099)
         );
  MUX2X1 U2243 ( .B(n2098), .A(n2095), .S(n21), .Y(n2102) );
  MUX2X1 U2244 ( .B(n2101), .A(n2086), .S(n23), .Y(n2235) );
  MUX2X1 U2245 ( .B(fifo_array[492]), .A(fifo_array[508]), .S(n2256), .Y(n2106) );
  MUX2X1 U2246 ( .B(fifo_array[460]), .A(fifo_array[476]), .S(n2256), .Y(n2105) );
  MUX2X1 U2247 ( .B(fifo_array[428]), .A(fifo_array[444]), .S(n2256), .Y(n2109) );
  MUX2X1 U2248 ( .B(fifo_array[396]), .A(fifo_array[412]), .S(n2256), .Y(n2108) );
  MUX2X1 U2249 ( .B(n2107), .A(n2104), .S(n21), .Y(n2118) );
  MUX2X1 U2250 ( .B(fifo_array[364]), .A(fifo_array[380]), .S(n2245), .Y(n2112) );
  MUX2X1 U2251 ( .B(fifo_array[332]), .A(fifo_array[348]), .S(n2242), .Y(n2111) );
  MUX2X1 U2252 ( .B(fifo_array[300]), .A(fifo_array[316]), .S(n2256), .Y(n2115) );
  MUX2X1 U2253 ( .B(fifo_array[268]), .A(fifo_array[284]), .S(n2244), .Y(n2114) );
  MUX2X1 U2254 ( .B(n2113), .A(n2110), .S(n21), .Y(n2117) );
  MUX2X1 U2255 ( .B(fifo_array[236]), .A(fifo_array[252]), .S(n2249), .Y(n2121) );
  MUX2X1 U2256 ( .B(fifo_array[204]), .A(fifo_array[220]), .S(n2252), .Y(n2120) );
  MUX2X1 U2257 ( .B(fifo_array[172]), .A(fifo_array[188]), .S(n2250), .Y(n2124) );
  MUX2X1 U2258 ( .B(fifo_array[140]), .A(fifo_array[156]), .S(n2251), .Y(n2123) );
  MUX2X1 U2259 ( .B(n2122), .A(n2119), .S(n21), .Y(n2133) );
  MUX2X1 U2260 ( .B(fifo_array[108]), .A(fifo_array[124]), .S(n2254), .Y(n2127) );
  MUX2X1 U2261 ( .B(fifo_array[76]), .A(fifo_array[92]), .S(n2241), .Y(n2126)
         );
  MUX2X1 U2262 ( .B(fifo_array[44]), .A(fifo_array[60]), .S(n2247), .Y(n2130)
         );
  MUX2X1 U2263 ( .B(fifo_array[12]), .A(fifo_array[28]), .S(n2248), .Y(n2129)
         );
  MUX2X1 U2264 ( .B(n2128), .A(n2125), .S(n21), .Y(n2132) );
  MUX2X1 U2265 ( .B(n2131), .A(n2116), .S(n23), .Y(n2236) );
  MUX2X1 U2266 ( .B(fifo_array[493]), .A(fifo_array[509]), .S(n2244), .Y(n2136) );
  MUX2X1 U2267 ( .B(fifo_array[461]), .A(fifo_array[477]), .S(n2255), .Y(n2135) );
  MUX2X1 U2268 ( .B(fifo_array[429]), .A(fifo_array[445]), .S(n2256), .Y(n2139) );
  MUX2X1 U2269 ( .B(fifo_array[397]), .A(fifo_array[413]), .S(n2242), .Y(n2138) );
  MUX2X1 U2270 ( .B(n2137), .A(n2134), .S(n21), .Y(n2148) );
  MUX2X1 U2271 ( .B(fifo_array[365]), .A(fifo_array[381]), .S(n2246), .Y(n2142) );
  MUX2X1 U2272 ( .B(fifo_array[333]), .A(fifo_array[349]), .S(n2243), .Y(n2141) );
  MUX2X1 U2273 ( .B(fifo_array[301]), .A(fifo_array[317]), .S(n2241), .Y(n2145) );
  MUX2X1 U2274 ( .B(fifo_array[269]), .A(fifo_array[285]), .S(n2245), .Y(n2144) );
  MUX2X1 U2275 ( .B(n2143), .A(n2140), .S(n21), .Y(n2147) );
  MUX2X1 U2276 ( .B(fifo_array[237]), .A(fifo_array[253]), .S(n2252), .Y(n2151) );
  MUX2X1 U2277 ( .B(fifo_array[205]), .A(fifo_array[221]), .S(n2253), .Y(n2150) );
  MUX2X1 U2278 ( .B(fifo_array[173]), .A(fifo_array[189]), .S(n2250), .Y(n2154) );
  MUX2X1 U2279 ( .B(fifo_array[141]), .A(fifo_array[157]), .S(n2253), .Y(n2153) );
  MUX2X1 U2280 ( .B(n2152), .A(n2149), .S(n21), .Y(n2163) );
  MUX2X1 U2281 ( .B(fifo_array[109]), .A(fifo_array[125]), .S(n2257), .Y(n2157) );
  MUX2X1 U2282 ( .B(fifo_array[77]), .A(fifo_array[93]), .S(n2257), .Y(n2156)
         );
  MUX2X1 U2283 ( .B(fifo_array[45]), .A(fifo_array[61]), .S(n2257), .Y(n2160)
         );
  MUX2X1 U2284 ( .B(fifo_array[13]), .A(fifo_array[29]), .S(n2257), .Y(n2159)
         );
  MUX2X1 U2285 ( .B(n2158), .A(n2155), .S(n21), .Y(n2162) );
  MUX2X1 U2286 ( .B(n2161), .A(n2146), .S(n23), .Y(n2237) );
  MUX2X1 U2287 ( .B(fifo_array[494]), .A(fifo_array[510]), .S(n2257), .Y(n2166) );
  MUX2X1 U2288 ( .B(fifo_array[462]), .A(fifo_array[478]), .S(n2257), .Y(n2165) );
  MUX2X1 U2289 ( .B(fifo_array[430]), .A(fifo_array[446]), .S(n2257), .Y(n2169) );
  MUX2X1 U2290 ( .B(fifo_array[398]), .A(fifo_array[414]), .S(n2257), .Y(n2168) );
  MUX2X1 U2291 ( .B(n2167), .A(n2164), .S(n21), .Y(n2178) );
  MUX2X1 U2292 ( .B(fifo_array[366]), .A(fifo_array[382]), .S(n2257), .Y(n2172) );
  MUX2X1 U2293 ( .B(fifo_array[334]), .A(fifo_array[350]), .S(n2257), .Y(n2171) );
  MUX2X1 U2294 ( .B(fifo_array[302]), .A(fifo_array[318]), .S(n2257), .Y(n2175) );
  MUX2X1 U2295 ( .B(fifo_array[270]), .A(fifo_array[286]), .S(n2257), .Y(n2174) );
  MUX2X1 U2296 ( .B(n2173), .A(n2170), .S(n21), .Y(n2177) );
  MUX2X1 U2297 ( .B(fifo_array[238]), .A(fifo_array[254]), .S(n2247), .Y(n2181) );
  MUX2X1 U2298 ( .B(fifo_array[206]), .A(fifo_array[222]), .S(n2249), .Y(n2180) );
  MUX2X1 U2299 ( .B(fifo_array[174]), .A(fifo_array[190]), .S(n2244), .Y(n2184) );
  MUX2X1 U2300 ( .B(fifo_array[142]), .A(fifo_array[158]), .S(n2243), .Y(n2183) );
  MUX2X1 U2301 ( .B(n2182), .A(n2179), .S(n21), .Y(n2193) );
  MUX2X1 U2302 ( .B(fifo_array[110]), .A(fifo_array[126]), .S(n2248), .Y(n2187) );
  MUX2X1 U2303 ( .B(fifo_array[78]), .A(fifo_array[94]), .S(n2243), .Y(n2186)
         );
  MUX2X1 U2304 ( .B(fifo_array[46]), .A(fifo_array[62]), .S(n2251), .Y(n2190)
         );
  MUX2X1 U2305 ( .B(fifo_array[14]), .A(fifo_array[30]), .S(n2254), .Y(n2189)
         );
  MUX2X1 U2306 ( .B(n2188), .A(n2185), .S(n21), .Y(n2192) );
  MUX2X1 U2307 ( .B(n2191), .A(n2176), .S(n23), .Y(n2238) );
  MUX2X1 U2308 ( .B(fifo_array[495]), .A(fifo_array[511]), .S(n2242), .Y(n2196) );
  MUX2X1 U2309 ( .B(fifo_array[463]), .A(fifo_array[479]), .S(n2245), .Y(n2195) );
  MUX2X1 U2310 ( .B(fifo_array[431]), .A(fifo_array[447]), .S(n2255), .Y(n2199) );
  MUX2X1 U2311 ( .B(fifo_array[399]), .A(fifo_array[415]), .S(n2246), .Y(n2198) );
  MUX2X1 U2312 ( .B(n2197), .A(n2194), .S(n21), .Y(n2208) );
  MUX2X1 U2313 ( .B(fifo_array[367]), .A(fifo_array[383]), .S(n2311), .Y(n2202) );
  MUX2X1 U2314 ( .B(fifo_array[335]), .A(fifo_array[351]), .S(n2257), .Y(n2201) );
  MUX2X1 U2315 ( .B(fifo_array[303]), .A(fifo_array[319]), .S(n2311), .Y(n2205) );
  MUX2X1 U2316 ( .B(fifo_array[271]), .A(fifo_array[287]), .S(n2311), .Y(n2204) );
  MUX2X1 U2317 ( .B(n2203), .A(n2200), .S(n21), .Y(n2207) );
  MUX2X1 U2318 ( .B(fifo_array[239]), .A(fifo_array[255]), .S(n2311), .Y(n2211) );
  MUX2X1 U2319 ( .B(fifo_array[207]), .A(fifo_array[223]), .S(n2311), .Y(n2210) );
  MUX2X1 U2320 ( .B(fifo_array[175]), .A(fifo_array[191]), .S(n2311), .Y(n2214) );
  MUX2X1 U2321 ( .B(fifo_array[143]), .A(fifo_array[159]), .S(n2311), .Y(n2213) );
  MUX2X1 U2322 ( .B(n2212), .A(n2209), .S(n21), .Y(n2223) );
  MUX2X1 U2323 ( .B(fifo_array[111]), .A(fifo_array[127]), .S(n2311), .Y(n2217) );
  MUX2X1 U2324 ( .B(fifo_array[79]), .A(fifo_array[95]), .S(n2311), .Y(n2216)
         );
  MUX2X1 U2325 ( .B(fifo_array[47]), .A(fifo_array[63]), .S(n2311), .Y(n2220)
         );
  MUX2X1 U2326 ( .B(fifo_array[15]), .A(fifo_array[31]), .S(n2311), .Y(n2219)
         );
  MUX2X1 U2327 ( .B(n2218), .A(n2215), .S(n21), .Y(n2222) );
  MUX2X1 U2328 ( .B(n2221), .A(n2206), .S(n23), .Y(n2239) );
  INVX1 U2329 ( .A(n2261), .Y(n2262) );
  XOR2X1 U2330 ( .A(r307_carry[4]), .B(wr_ptr[4]), .Y(n53) );
  XOR2X1 U2331 ( .A(r308_carry[4]), .B(n23), .Y(n58) );
  XOR2X1 U2332 ( .A(add_45_carry[5]), .B(fillcount[5]), .Y(n70) );
  OAI21X1 U2333 ( .A(n77), .B(n2350), .C(n1708), .Y(n78) );
  OAI21X1 U2334 ( .A(n2313), .B(n2318), .C(n1666), .Y(n79) );
  OAI21X1 U2335 ( .A(n2314), .B(n2317), .C(n1709), .Y(n80) );
  XNOR2X1 U2336 ( .A(fillcount[4]), .B(n1709), .Y(n81) );
  XNOR2X1 U2337 ( .A(fillcount[5]), .B(n2316), .Y(n82) );
endmodule


module FIFO_DEPTH_P25_WIDTH34 ( clk, reset, data_in, put, get, data_out, empty, 
        full, fillcount );
  input [33:0] data_in;
  output [33:0] data_out;
  output [5:0] fillcount;
  input clk, reset, put, get;
  output empty, full;
  wire   n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n68, n69, n70,
         n71, n73, n74, n75, n76, n84, n85, n86, n87, n88, n95, n96, n97, n98,
         n99, n100, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n72, n77, n78, n79, n80, n81, n82, n83, n89, n90, n91,
         n92, n93, n94, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n1304, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814;
  wire   [4:0] wr_ptr;
  wire   [1087:0] fifo_array;
  wire   [5:2] add_45_carry;
  wire   [4:2] r308_carry;
  wire   [4:2] r307_carry;

  DFFPOSX1 full_reg ( .D(n2463), .CLK(clk), .Q(full) );
  DFFPOSX1 fillcount_reg_5_ ( .D(n2462), .CLK(clk), .Q(fillcount[5]) );
  DFFPOSX1 empty_reg ( .D(n2461), .CLK(clk), .Q(empty) );
  DFFPOSX1 wr_ptr_reg_0_ ( .D(n2455), .CLK(clk), .Q(wr_ptr[0]) );
  DFFPOSX1 wr_ptr_reg_1_ ( .D(n2454), .CLK(clk), .Q(wr_ptr[1]) );
  DFFPOSX1 wr_ptr_reg_2_ ( .D(n2453), .CLK(clk), .Q(wr_ptr[2]) );
  DFFPOSX1 wr_ptr_reg_3_ ( .D(n2452), .CLK(clk), .Q(wr_ptr[3]) );
  DFFPOSX1 wr_ptr_reg_4_ ( .D(n2451), .CLK(clk), .Q(wr_ptr[4]) );
  DFFPOSX1 data_out_reg_0_ ( .D(n4766), .CLK(clk), .Q(data_out[0]) );
  DFFPOSX1 data_out_reg_1_ ( .D(n4767), .CLK(clk), .Q(data_out[1]) );
  DFFPOSX1 data_out_reg_2_ ( .D(n4768), .CLK(clk), .Q(data_out[2]) );
  DFFPOSX1 data_out_reg_3_ ( .D(n4769), .CLK(clk), .Q(data_out[3]) );
  DFFPOSX1 data_out_reg_4_ ( .D(n4770), .CLK(clk), .Q(data_out[4]) );
  DFFPOSX1 data_out_reg_5_ ( .D(n4771), .CLK(clk), .Q(data_out[5]) );
  DFFPOSX1 data_out_reg_6_ ( .D(n4772), .CLK(clk), .Q(data_out[6]) );
  DFFPOSX1 data_out_reg_7_ ( .D(n4773), .CLK(clk), .Q(data_out[7]) );
  DFFPOSX1 data_out_reg_8_ ( .D(n4774), .CLK(clk), .Q(data_out[8]) );
  DFFPOSX1 data_out_reg_9_ ( .D(n4775), .CLK(clk), .Q(data_out[9]) );
  DFFPOSX1 data_out_reg_10_ ( .D(n4776), .CLK(clk), .Q(data_out[10]) );
  DFFPOSX1 data_out_reg_11_ ( .D(n4777), .CLK(clk), .Q(data_out[11]) );
  DFFPOSX1 data_out_reg_12_ ( .D(n4778), .CLK(clk), .Q(data_out[12]) );
  DFFPOSX1 data_out_reg_13_ ( .D(n4779), .CLK(clk), .Q(data_out[13]) );
  DFFPOSX1 data_out_reg_14_ ( .D(n4780), .CLK(clk), .Q(data_out[14]) );
  DFFPOSX1 data_out_reg_15_ ( .D(n4781), .CLK(clk), .Q(data_out[15]) );
  DFFPOSX1 data_out_reg_16_ ( .D(n4782), .CLK(clk), .Q(data_out[16]) );
  DFFPOSX1 data_out_reg_17_ ( .D(n4783), .CLK(clk), .Q(data_out[17]) );
  DFFPOSX1 data_out_reg_18_ ( .D(n4784), .CLK(clk), .Q(data_out[18]) );
  DFFPOSX1 data_out_reg_19_ ( .D(n4785), .CLK(clk), .Q(data_out[19]) );
  DFFPOSX1 data_out_reg_20_ ( .D(n4786), .CLK(clk), .Q(data_out[20]) );
  DFFPOSX1 data_out_reg_21_ ( .D(n4787), .CLK(clk), .Q(data_out[21]) );
  DFFPOSX1 data_out_reg_22_ ( .D(n4788), .CLK(clk), .Q(data_out[22]) );
  DFFPOSX1 data_out_reg_23_ ( .D(n4789), .CLK(clk), .Q(data_out[23]) );
  DFFPOSX1 data_out_reg_24_ ( .D(n4790), .CLK(clk), .Q(data_out[24]) );
  DFFPOSX1 data_out_reg_25_ ( .D(n4791), .CLK(clk), .Q(data_out[25]) );
  DFFPOSX1 data_out_reg_26_ ( .D(n4792), .CLK(clk), .Q(data_out[26]) );
  DFFPOSX1 data_out_reg_27_ ( .D(n4793), .CLK(clk), .Q(data_out[27]) );
  DFFPOSX1 data_out_reg_28_ ( .D(n4794), .CLK(clk), .Q(data_out[28]) );
  DFFPOSX1 data_out_reg_29_ ( .D(n4795), .CLK(clk), .Q(data_out[29]) );
  DFFPOSX1 data_out_reg_30_ ( .D(n4796), .CLK(clk), .Q(data_out[30]) );
  DFFPOSX1 data_out_reg_31_ ( .D(n4797), .CLK(clk), .Q(data_out[31]) );
  DFFPOSX1 data_out_reg_32_ ( .D(n4798), .CLK(clk), .Q(data_out[32]) );
  DFFPOSX1 data_out_reg_33_ ( .D(n4799), .CLK(clk), .Q(data_out[33]) );
  DFFPOSX1 rd_ptr_reg_0_ ( .D(n4800), .CLK(clk), .Q(n19) );
  DFFPOSX1 rd_ptr_reg_1_ ( .D(n4801), .CLK(clk), .Q(n20) );
  DFFPOSX1 rd_ptr_reg_2_ ( .D(n4802), .CLK(clk), .Q(n21) );
  DFFPOSX1 rd_ptr_reg_3_ ( .D(n4803), .CLK(clk), .Q(n22) );
  DFFPOSX1 rd_ptr_reg_4_ ( .D(n4804), .CLK(clk), .Q(n23) );
  DFFPOSX1 fillcount_reg_0_ ( .D(n2460), .CLK(clk), .Q(fillcount[0]) );
  DFFPOSX1 fillcount_reg_4_ ( .D(n2456), .CLK(clk), .Q(fillcount[4]) );
  DFFPOSX1 fillcount_reg_1_ ( .D(n2459), .CLK(clk), .Q(fillcount[1]) );
  DFFPOSX1 fillcount_reg_2_ ( .D(n2458), .CLK(clk), .Q(fillcount[2]) );
  DFFPOSX1 fillcount_reg_3_ ( .D(n2457), .CLK(clk), .Q(fillcount[3]) );
  DFFPOSX1 fifo_array_reg_31__33_ ( .D(n2450), .CLK(clk), .Q(fifo_array[1087])
         );
  DFFPOSX1 fifo_array_reg_31__32_ ( .D(n2449), .CLK(clk), .Q(fifo_array[1086])
         );
  DFFPOSX1 fifo_array_reg_31__31_ ( .D(n2448), .CLK(clk), .Q(fifo_array[1085])
         );
  DFFPOSX1 fifo_array_reg_31__30_ ( .D(n2447), .CLK(clk), .Q(fifo_array[1084])
         );
  DFFPOSX1 fifo_array_reg_31__29_ ( .D(n2446), .CLK(clk), .Q(fifo_array[1083])
         );
  DFFPOSX1 fifo_array_reg_31__28_ ( .D(n2445), .CLK(clk), .Q(fifo_array[1082])
         );
  DFFPOSX1 fifo_array_reg_31__27_ ( .D(n2444), .CLK(clk), .Q(fifo_array[1081])
         );
  DFFPOSX1 fifo_array_reg_31__26_ ( .D(n2443), .CLK(clk), .Q(fifo_array[1080])
         );
  DFFPOSX1 fifo_array_reg_31__25_ ( .D(n2442), .CLK(clk), .Q(fifo_array[1079])
         );
  DFFPOSX1 fifo_array_reg_31__24_ ( .D(n2441), .CLK(clk), .Q(fifo_array[1078])
         );
  DFFPOSX1 fifo_array_reg_31__23_ ( .D(n2440), .CLK(clk), .Q(fifo_array[1077])
         );
  DFFPOSX1 fifo_array_reg_31__22_ ( .D(n2439), .CLK(clk), .Q(fifo_array[1076])
         );
  DFFPOSX1 fifo_array_reg_31__21_ ( .D(n2438), .CLK(clk), .Q(fifo_array[1075])
         );
  DFFPOSX1 fifo_array_reg_31__20_ ( .D(n2437), .CLK(clk), .Q(fifo_array[1074])
         );
  DFFPOSX1 fifo_array_reg_31__19_ ( .D(n2436), .CLK(clk), .Q(fifo_array[1073])
         );
  DFFPOSX1 fifo_array_reg_31__18_ ( .D(n2435), .CLK(clk), .Q(fifo_array[1072])
         );
  DFFPOSX1 fifo_array_reg_31__17_ ( .D(n2434), .CLK(clk), .Q(fifo_array[1071])
         );
  DFFPOSX1 fifo_array_reg_31__16_ ( .D(n2433), .CLK(clk), .Q(fifo_array[1070])
         );
  DFFPOSX1 fifo_array_reg_31__15_ ( .D(n2432), .CLK(clk), .Q(fifo_array[1069])
         );
  DFFPOSX1 fifo_array_reg_31__14_ ( .D(n2431), .CLK(clk), .Q(fifo_array[1068])
         );
  DFFPOSX1 fifo_array_reg_31__13_ ( .D(n2430), .CLK(clk), .Q(fifo_array[1067])
         );
  DFFPOSX1 fifo_array_reg_31__12_ ( .D(n2429), .CLK(clk), .Q(fifo_array[1066])
         );
  DFFPOSX1 fifo_array_reg_31__11_ ( .D(n2428), .CLK(clk), .Q(fifo_array[1065])
         );
  DFFPOSX1 fifo_array_reg_31__10_ ( .D(n2427), .CLK(clk), .Q(fifo_array[1064])
         );
  DFFPOSX1 fifo_array_reg_31__9_ ( .D(n2426), .CLK(clk), .Q(fifo_array[1063])
         );
  DFFPOSX1 fifo_array_reg_31__8_ ( .D(n2425), .CLK(clk), .Q(fifo_array[1062])
         );
  DFFPOSX1 fifo_array_reg_31__7_ ( .D(n2424), .CLK(clk), .Q(fifo_array[1061])
         );
  DFFPOSX1 fifo_array_reg_31__6_ ( .D(n2423), .CLK(clk), .Q(fifo_array[1060])
         );
  DFFPOSX1 fifo_array_reg_31__5_ ( .D(n2422), .CLK(clk), .Q(fifo_array[1059])
         );
  DFFPOSX1 fifo_array_reg_31__4_ ( .D(n2421), .CLK(clk), .Q(fifo_array[1058])
         );
  DFFPOSX1 fifo_array_reg_31__3_ ( .D(n2420), .CLK(clk), .Q(fifo_array[1057])
         );
  DFFPOSX1 fifo_array_reg_31__2_ ( .D(n2419), .CLK(clk), .Q(fifo_array[1056])
         );
  DFFPOSX1 fifo_array_reg_31__1_ ( .D(n2418), .CLK(clk), .Q(fifo_array[1055])
         );
  DFFPOSX1 fifo_array_reg_31__0_ ( .D(n2417), .CLK(clk), .Q(fifo_array[1054])
         );
  DFFPOSX1 fifo_array_reg_30__33_ ( .D(n2416), .CLK(clk), .Q(fifo_array[1053])
         );
  DFFPOSX1 fifo_array_reg_30__32_ ( .D(n2415), .CLK(clk), .Q(fifo_array[1052])
         );
  DFFPOSX1 fifo_array_reg_30__31_ ( .D(n2414), .CLK(clk), .Q(fifo_array[1051])
         );
  DFFPOSX1 fifo_array_reg_30__30_ ( .D(n2413), .CLK(clk), .Q(fifo_array[1050])
         );
  DFFPOSX1 fifo_array_reg_30__29_ ( .D(n2412), .CLK(clk), .Q(fifo_array[1049])
         );
  DFFPOSX1 fifo_array_reg_30__28_ ( .D(n2411), .CLK(clk), .Q(fifo_array[1048])
         );
  DFFPOSX1 fifo_array_reg_30__27_ ( .D(n2410), .CLK(clk), .Q(fifo_array[1047])
         );
  DFFPOSX1 fifo_array_reg_30__26_ ( .D(n2409), .CLK(clk), .Q(fifo_array[1046])
         );
  DFFPOSX1 fifo_array_reg_30__25_ ( .D(n2408), .CLK(clk), .Q(fifo_array[1045])
         );
  DFFPOSX1 fifo_array_reg_30__24_ ( .D(n2407), .CLK(clk), .Q(fifo_array[1044])
         );
  DFFPOSX1 fifo_array_reg_30__23_ ( .D(n2406), .CLK(clk), .Q(fifo_array[1043])
         );
  DFFPOSX1 fifo_array_reg_30__22_ ( .D(n2405), .CLK(clk), .Q(fifo_array[1042])
         );
  DFFPOSX1 fifo_array_reg_30__21_ ( .D(n2404), .CLK(clk), .Q(fifo_array[1041])
         );
  DFFPOSX1 fifo_array_reg_30__20_ ( .D(n2403), .CLK(clk), .Q(fifo_array[1040])
         );
  DFFPOSX1 fifo_array_reg_30__19_ ( .D(n2402), .CLK(clk), .Q(fifo_array[1039])
         );
  DFFPOSX1 fifo_array_reg_30__18_ ( .D(n2401), .CLK(clk), .Q(fifo_array[1038])
         );
  DFFPOSX1 fifo_array_reg_30__17_ ( .D(n2400), .CLK(clk), .Q(fifo_array[1037])
         );
  DFFPOSX1 fifo_array_reg_30__16_ ( .D(n2399), .CLK(clk), .Q(fifo_array[1036])
         );
  DFFPOSX1 fifo_array_reg_30__15_ ( .D(n2398), .CLK(clk), .Q(fifo_array[1035])
         );
  DFFPOSX1 fifo_array_reg_30__14_ ( .D(n2397), .CLK(clk), .Q(fifo_array[1034])
         );
  DFFPOSX1 fifo_array_reg_30__13_ ( .D(n2396), .CLK(clk), .Q(fifo_array[1033])
         );
  DFFPOSX1 fifo_array_reg_30__12_ ( .D(n2395), .CLK(clk), .Q(fifo_array[1032])
         );
  DFFPOSX1 fifo_array_reg_30__11_ ( .D(n2394), .CLK(clk), .Q(fifo_array[1031])
         );
  DFFPOSX1 fifo_array_reg_30__10_ ( .D(n2393), .CLK(clk), .Q(fifo_array[1030])
         );
  DFFPOSX1 fifo_array_reg_30__9_ ( .D(n2392), .CLK(clk), .Q(fifo_array[1029])
         );
  DFFPOSX1 fifo_array_reg_30__8_ ( .D(n2391), .CLK(clk), .Q(fifo_array[1028])
         );
  DFFPOSX1 fifo_array_reg_30__7_ ( .D(n2390), .CLK(clk), .Q(fifo_array[1027])
         );
  DFFPOSX1 fifo_array_reg_30__6_ ( .D(n2389), .CLK(clk), .Q(fifo_array[1026])
         );
  DFFPOSX1 fifo_array_reg_30__5_ ( .D(n2388), .CLK(clk), .Q(fifo_array[1025])
         );
  DFFPOSX1 fifo_array_reg_30__4_ ( .D(n2387), .CLK(clk), .Q(fifo_array[1024])
         );
  DFFPOSX1 fifo_array_reg_30__3_ ( .D(n2386), .CLK(clk), .Q(fifo_array[1023])
         );
  DFFPOSX1 fifo_array_reg_30__2_ ( .D(n2385), .CLK(clk), .Q(fifo_array[1022])
         );
  DFFPOSX1 fifo_array_reg_30__1_ ( .D(n2384), .CLK(clk), .Q(fifo_array[1021])
         );
  DFFPOSX1 fifo_array_reg_30__0_ ( .D(n2383), .CLK(clk), .Q(fifo_array[1020])
         );
  DFFPOSX1 fifo_array_reg_29__33_ ( .D(n2382), .CLK(clk), .Q(fifo_array[1019])
         );
  DFFPOSX1 fifo_array_reg_29__32_ ( .D(n2381), .CLK(clk), .Q(fifo_array[1018])
         );
  DFFPOSX1 fifo_array_reg_29__31_ ( .D(n2380), .CLK(clk), .Q(fifo_array[1017])
         );
  DFFPOSX1 fifo_array_reg_29__30_ ( .D(n2379), .CLK(clk), .Q(fifo_array[1016])
         );
  DFFPOSX1 fifo_array_reg_29__29_ ( .D(n2378), .CLK(clk), .Q(fifo_array[1015])
         );
  DFFPOSX1 fifo_array_reg_29__28_ ( .D(n2377), .CLK(clk), .Q(fifo_array[1014])
         );
  DFFPOSX1 fifo_array_reg_29__27_ ( .D(n2376), .CLK(clk), .Q(fifo_array[1013])
         );
  DFFPOSX1 fifo_array_reg_29__26_ ( .D(n2375), .CLK(clk), .Q(fifo_array[1012])
         );
  DFFPOSX1 fifo_array_reg_29__25_ ( .D(n2374), .CLK(clk), .Q(fifo_array[1011])
         );
  DFFPOSX1 fifo_array_reg_29__24_ ( .D(n2373), .CLK(clk), .Q(fifo_array[1010])
         );
  DFFPOSX1 fifo_array_reg_29__23_ ( .D(n2372), .CLK(clk), .Q(fifo_array[1009])
         );
  DFFPOSX1 fifo_array_reg_29__22_ ( .D(n2371), .CLK(clk), .Q(fifo_array[1008])
         );
  DFFPOSX1 fifo_array_reg_29__21_ ( .D(n2370), .CLK(clk), .Q(fifo_array[1007])
         );
  DFFPOSX1 fifo_array_reg_29__20_ ( .D(n2369), .CLK(clk), .Q(fifo_array[1006])
         );
  DFFPOSX1 fifo_array_reg_29__19_ ( .D(n2368), .CLK(clk), .Q(fifo_array[1005])
         );
  DFFPOSX1 fifo_array_reg_29__18_ ( .D(n2367), .CLK(clk), .Q(fifo_array[1004])
         );
  DFFPOSX1 fifo_array_reg_29__17_ ( .D(n2366), .CLK(clk), .Q(fifo_array[1003])
         );
  DFFPOSX1 fifo_array_reg_29__16_ ( .D(n2365), .CLK(clk), .Q(fifo_array[1002])
         );
  DFFPOSX1 fifo_array_reg_29__15_ ( .D(n2364), .CLK(clk), .Q(fifo_array[1001])
         );
  DFFPOSX1 fifo_array_reg_29__14_ ( .D(n2363), .CLK(clk), .Q(fifo_array[1000])
         );
  DFFPOSX1 fifo_array_reg_29__13_ ( .D(n2362), .CLK(clk), .Q(fifo_array[999])
         );
  DFFPOSX1 fifo_array_reg_29__12_ ( .D(n2361), .CLK(clk), .Q(fifo_array[998])
         );
  DFFPOSX1 fifo_array_reg_29__11_ ( .D(n2360), .CLK(clk), .Q(fifo_array[997])
         );
  DFFPOSX1 fifo_array_reg_29__10_ ( .D(n2359), .CLK(clk), .Q(fifo_array[996])
         );
  DFFPOSX1 fifo_array_reg_29__9_ ( .D(n2358), .CLK(clk), .Q(fifo_array[995])
         );
  DFFPOSX1 fifo_array_reg_29__8_ ( .D(n2357), .CLK(clk), .Q(fifo_array[994])
         );
  DFFPOSX1 fifo_array_reg_29__7_ ( .D(n2356), .CLK(clk), .Q(fifo_array[993])
         );
  DFFPOSX1 fifo_array_reg_29__6_ ( .D(n2355), .CLK(clk), .Q(fifo_array[992])
         );
  DFFPOSX1 fifo_array_reg_29__5_ ( .D(n2354), .CLK(clk), .Q(fifo_array[991])
         );
  DFFPOSX1 fifo_array_reg_29__4_ ( .D(n2353), .CLK(clk), .Q(fifo_array[990])
         );
  DFFPOSX1 fifo_array_reg_29__3_ ( .D(n2352), .CLK(clk), .Q(fifo_array[989])
         );
  DFFPOSX1 fifo_array_reg_29__2_ ( .D(n2351), .CLK(clk), .Q(fifo_array[988])
         );
  DFFPOSX1 fifo_array_reg_29__1_ ( .D(n2350), .CLK(clk), .Q(fifo_array[987])
         );
  DFFPOSX1 fifo_array_reg_29__0_ ( .D(n2349), .CLK(clk), .Q(fifo_array[986])
         );
  DFFPOSX1 fifo_array_reg_28__33_ ( .D(n2348), .CLK(clk), .Q(fifo_array[985])
         );
  DFFPOSX1 fifo_array_reg_28__32_ ( .D(n2347), .CLK(clk), .Q(fifo_array[984])
         );
  DFFPOSX1 fifo_array_reg_28__31_ ( .D(n2346), .CLK(clk), .Q(fifo_array[983])
         );
  DFFPOSX1 fifo_array_reg_28__30_ ( .D(n2345), .CLK(clk), .Q(fifo_array[982])
         );
  DFFPOSX1 fifo_array_reg_28__29_ ( .D(n2344), .CLK(clk), .Q(fifo_array[981])
         );
  DFFPOSX1 fifo_array_reg_28__28_ ( .D(n2343), .CLK(clk), .Q(fifo_array[980])
         );
  DFFPOSX1 fifo_array_reg_28__27_ ( .D(n2342), .CLK(clk), .Q(fifo_array[979])
         );
  DFFPOSX1 fifo_array_reg_28__26_ ( .D(n2341), .CLK(clk), .Q(fifo_array[978])
         );
  DFFPOSX1 fifo_array_reg_28__25_ ( .D(n2340), .CLK(clk), .Q(fifo_array[977])
         );
  DFFPOSX1 fifo_array_reg_28__24_ ( .D(n2339), .CLK(clk), .Q(fifo_array[976])
         );
  DFFPOSX1 fifo_array_reg_28__23_ ( .D(n2338), .CLK(clk), .Q(fifo_array[975])
         );
  DFFPOSX1 fifo_array_reg_28__22_ ( .D(n2337), .CLK(clk), .Q(fifo_array[974])
         );
  DFFPOSX1 fifo_array_reg_28__21_ ( .D(n2336), .CLK(clk), .Q(fifo_array[973])
         );
  DFFPOSX1 fifo_array_reg_28__20_ ( .D(n2335), .CLK(clk), .Q(fifo_array[972])
         );
  DFFPOSX1 fifo_array_reg_28__19_ ( .D(n2334), .CLK(clk), .Q(fifo_array[971])
         );
  DFFPOSX1 fifo_array_reg_28__18_ ( .D(n2333), .CLK(clk), .Q(fifo_array[970])
         );
  DFFPOSX1 fifo_array_reg_28__17_ ( .D(n2332), .CLK(clk), .Q(fifo_array[969])
         );
  DFFPOSX1 fifo_array_reg_28__16_ ( .D(n2331), .CLK(clk), .Q(fifo_array[968])
         );
  DFFPOSX1 fifo_array_reg_28__15_ ( .D(n2330), .CLK(clk), .Q(fifo_array[967])
         );
  DFFPOSX1 fifo_array_reg_28__14_ ( .D(n2329), .CLK(clk), .Q(fifo_array[966])
         );
  DFFPOSX1 fifo_array_reg_28__13_ ( .D(n2328), .CLK(clk), .Q(fifo_array[965])
         );
  DFFPOSX1 fifo_array_reg_28__12_ ( .D(n2327), .CLK(clk), .Q(fifo_array[964])
         );
  DFFPOSX1 fifo_array_reg_28__11_ ( .D(n2326), .CLK(clk), .Q(fifo_array[963])
         );
  DFFPOSX1 fifo_array_reg_28__10_ ( .D(n2325), .CLK(clk), .Q(fifo_array[962])
         );
  DFFPOSX1 fifo_array_reg_28__9_ ( .D(n2324), .CLK(clk), .Q(fifo_array[961])
         );
  DFFPOSX1 fifo_array_reg_28__8_ ( .D(n2323), .CLK(clk), .Q(fifo_array[960])
         );
  DFFPOSX1 fifo_array_reg_28__7_ ( .D(n2322), .CLK(clk), .Q(fifo_array[959])
         );
  DFFPOSX1 fifo_array_reg_28__6_ ( .D(n2321), .CLK(clk), .Q(fifo_array[958])
         );
  DFFPOSX1 fifo_array_reg_28__5_ ( .D(n2320), .CLK(clk), .Q(fifo_array[957])
         );
  DFFPOSX1 fifo_array_reg_28__4_ ( .D(n2319), .CLK(clk), .Q(fifo_array[956])
         );
  DFFPOSX1 fifo_array_reg_28__3_ ( .D(n2318), .CLK(clk), .Q(fifo_array[955])
         );
  DFFPOSX1 fifo_array_reg_28__2_ ( .D(n2317), .CLK(clk), .Q(fifo_array[954])
         );
  DFFPOSX1 fifo_array_reg_28__1_ ( .D(n2316), .CLK(clk), .Q(fifo_array[953])
         );
  DFFPOSX1 fifo_array_reg_28__0_ ( .D(n2315), .CLK(clk), .Q(fifo_array[952])
         );
  DFFPOSX1 fifo_array_reg_27__33_ ( .D(n2314), .CLK(clk), .Q(fifo_array[951])
         );
  DFFPOSX1 fifo_array_reg_27__32_ ( .D(n2313), .CLK(clk), .Q(fifo_array[950])
         );
  DFFPOSX1 fifo_array_reg_27__31_ ( .D(n2312), .CLK(clk), .Q(fifo_array[949])
         );
  DFFPOSX1 fifo_array_reg_27__30_ ( .D(n2311), .CLK(clk), .Q(fifo_array[948])
         );
  DFFPOSX1 fifo_array_reg_27__29_ ( .D(n2310), .CLK(clk), .Q(fifo_array[947])
         );
  DFFPOSX1 fifo_array_reg_27__28_ ( .D(n2309), .CLK(clk), .Q(fifo_array[946])
         );
  DFFPOSX1 fifo_array_reg_27__27_ ( .D(n2308), .CLK(clk), .Q(fifo_array[945])
         );
  DFFPOSX1 fifo_array_reg_27__26_ ( .D(n2307), .CLK(clk), .Q(fifo_array[944])
         );
  DFFPOSX1 fifo_array_reg_27__25_ ( .D(n2306), .CLK(clk), .Q(fifo_array[943])
         );
  DFFPOSX1 fifo_array_reg_27__24_ ( .D(n2305), .CLK(clk), .Q(fifo_array[942])
         );
  DFFPOSX1 fifo_array_reg_27__23_ ( .D(n2304), .CLK(clk), .Q(fifo_array[941])
         );
  DFFPOSX1 fifo_array_reg_27__22_ ( .D(n2303), .CLK(clk), .Q(fifo_array[940])
         );
  DFFPOSX1 fifo_array_reg_27__21_ ( .D(n2302), .CLK(clk), .Q(fifo_array[939])
         );
  DFFPOSX1 fifo_array_reg_27__20_ ( .D(n2301), .CLK(clk), .Q(fifo_array[938])
         );
  DFFPOSX1 fifo_array_reg_27__19_ ( .D(n2300), .CLK(clk), .Q(fifo_array[937])
         );
  DFFPOSX1 fifo_array_reg_27__18_ ( .D(n2299), .CLK(clk), .Q(fifo_array[936])
         );
  DFFPOSX1 fifo_array_reg_27__17_ ( .D(n2298), .CLK(clk), .Q(fifo_array[935])
         );
  DFFPOSX1 fifo_array_reg_27__16_ ( .D(n2297), .CLK(clk), .Q(fifo_array[934])
         );
  DFFPOSX1 fifo_array_reg_27__15_ ( .D(n2296), .CLK(clk), .Q(fifo_array[933])
         );
  DFFPOSX1 fifo_array_reg_27__14_ ( .D(n2295), .CLK(clk), .Q(fifo_array[932])
         );
  DFFPOSX1 fifo_array_reg_27__13_ ( .D(n2294), .CLK(clk), .Q(fifo_array[931])
         );
  DFFPOSX1 fifo_array_reg_27__12_ ( .D(n2293), .CLK(clk), .Q(fifo_array[930])
         );
  DFFPOSX1 fifo_array_reg_27__11_ ( .D(n2292), .CLK(clk), .Q(fifo_array[929])
         );
  DFFPOSX1 fifo_array_reg_27__10_ ( .D(n2291), .CLK(clk), .Q(fifo_array[928])
         );
  DFFPOSX1 fifo_array_reg_27__9_ ( .D(n2290), .CLK(clk), .Q(fifo_array[927])
         );
  DFFPOSX1 fifo_array_reg_27__8_ ( .D(n2289), .CLK(clk), .Q(fifo_array[926])
         );
  DFFPOSX1 fifo_array_reg_27__7_ ( .D(n2288), .CLK(clk), .Q(fifo_array[925])
         );
  DFFPOSX1 fifo_array_reg_27__6_ ( .D(n2287), .CLK(clk), .Q(fifo_array[924])
         );
  DFFPOSX1 fifo_array_reg_27__5_ ( .D(n2286), .CLK(clk), .Q(fifo_array[923])
         );
  DFFPOSX1 fifo_array_reg_27__4_ ( .D(n2285), .CLK(clk), .Q(fifo_array[922])
         );
  DFFPOSX1 fifo_array_reg_27__3_ ( .D(n2284), .CLK(clk), .Q(fifo_array[921])
         );
  DFFPOSX1 fifo_array_reg_27__2_ ( .D(n2283), .CLK(clk), .Q(fifo_array[920])
         );
  DFFPOSX1 fifo_array_reg_27__1_ ( .D(n2282), .CLK(clk), .Q(fifo_array[919])
         );
  DFFPOSX1 fifo_array_reg_27__0_ ( .D(n2281), .CLK(clk), .Q(fifo_array[918])
         );
  DFFPOSX1 fifo_array_reg_26__33_ ( .D(n2280), .CLK(clk), .Q(fifo_array[917])
         );
  DFFPOSX1 fifo_array_reg_26__32_ ( .D(n2279), .CLK(clk), .Q(fifo_array[916])
         );
  DFFPOSX1 fifo_array_reg_26__31_ ( .D(n2278), .CLK(clk), .Q(fifo_array[915])
         );
  DFFPOSX1 fifo_array_reg_26__30_ ( .D(n2277), .CLK(clk), .Q(fifo_array[914])
         );
  DFFPOSX1 fifo_array_reg_26__29_ ( .D(n2276), .CLK(clk), .Q(fifo_array[913])
         );
  DFFPOSX1 fifo_array_reg_26__28_ ( .D(n2275), .CLK(clk), .Q(fifo_array[912])
         );
  DFFPOSX1 fifo_array_reg_26__27_ ( .D(n2274), .CLK(clk), .Q(fifo_array[911])
         );
  DFFPOSX1 fifo_array_reg_26__26_ ( .D(n2273), .CLK(clk), .Q(fifo_array[910])
         );
  DFFPOSX1 fifo_array_reg_26__25_ ( .D(n2272), .CLK(clk), .Q(fifo_array[909])
         );
  DFFPOSX1 fifo_array_reg_26__24_ ( .D(n2271), .CLK(clk), .Q(fifo_array[908])
         );
  DFFPOSX1 fifo_array_reg_26__23_ ( .D(n2270), .CLK(clk), .Q(fifo_array[907])
         );
  DFFPOSX1 fifo_array_reg_26__22_ ( .D(n2269), .CLK(clk), .Q(fifo_array[906])
         );
  DFFPOSX1 fifo_array_reg_26__21_ ( .D(n2268), .CLK(clk), .Q(fifo_array[905])
         );
  DFFPOSX1 fifo_array_reg_26__20_ ( .D(n2267), .CLK(clk), .Q(fifo_array[904])
         );
  DFFPOSX1 fifo_array_reg_26__19_ ( .D(n2266), .CLK(clk), .Q(fifo_array[903])
         );
  DFFPOSX1 fifo_array_reg_26__18_ ( .D(n2265), .CLK(clk), .Q(fifo_array[902])
         );
  DFFPOSX1 fifo_array_reg_26__17_ ( .D(n2264), .CLK(clk), .Q(fifo_array[901])
         );
  DFFPOSX1 fifo_array_reg_26__16_ ( .D(n2263), .CLK(clk), .Q(fifo_array[900])
         );
  DFFPOSX1 fifo_array_reg_26__15_ ( .D(n2262), .CLK(clk), .Q(fifo_array[899])
         );
  DFFPOSX1 fifo_array_reg_26__14_ ( .D(n2261), .CLK(clk), .Q(fifo_array[898])
         );
  DFFPOSX1 fifo_array_reg_26__13_ ( .D(n2260), .CLK(clk), .Q(fifo_array[897])
         );
  DFFPOSX1 fifo_array_reg_26__12_ ( .D(n2259), .CLK(clk), .Q(fifo_array[896])
         );
  DFFPOSX1 fifo_array_reg_26__11_ ( .D(n2258), .CLK(clk), .Q(fifo_array[895])
         );
  DFFPOSX1 fifo_array_reg_26__10_ ( .D(n2257), .CLK(clk), .Q(fifo_array[894])
         );
  DFFPOSX1 fifo_array_reg_26__9_ ( .D(n2256), .CLK(clk), .Q(fifo_array[893])
         );
  DFFPOSX1 fifo_array_reg_26__8_ ( .D(n2255), .CLK(clk), .Q(fifo_array[892])
         );
  DFFPOSX1 fifo_array_reg_26__7_ ( .D(n2254), .CLK(clk), .Q(fifo_array[891])
         );
  DFFPOSX1 fifo_array_reg_26__6_ ( .D(n2253), .CLK(clk), .Q(fifo_array[890])
         );
  DFFPOSX1 fifo_array_reg_26__5_ ( .D(n2252), .CLK(clk), .Q(fifo_array[889])
         );
  DFFPOSX1 fifo_array_reg_26__4_ ( .D(n2251), .CLK(clk), .Q(fifo_array[888])
         );
  DFFPOSX1 fifo_array_reg_26__3_ ( .D(n2250), .CLK(clk), .Q(fifo_array[887])
         );
  DFFPOSX1 fifo_array_reg_26__2_ ( .D(n2249), .CLK(clk), .Q(fifo_array[886])
         );
  DFFPOSX1 fifo_array_reg_26__1_ ( .D(n2248), .CLK(clk), .Q(fifo_array[885])
         );
  DFFPOSX1 fifo_array_reg_26__0_ ( .D(n2247), .CLK(clk), .Q(fifo_array[884])
         );
  DFFPOSX1 fifo_array_reg_25__33_ ( .D(n2246), .CLK(clk), .Q(fifo_array[883])
         );
  DFFPOSX1 fifo_array_reg_25__32_ ( .D(n2245), .CLK(clk), .Q(fifo_array[882])
         );
  DFFPOSX1 fifo_array_reg_25__31_ ( .D(n2244), .CLK(clk), .Q(fifo_array[881])
         );
  DFFPOSX1 fifo_array_reg_25__30_ ( .D(n2243), .CLK(clk), .Q(fifo_array[880])
         );
  DFFPOSX1 fifo_array_reg_25__29_ ( .D(n2242), .CLK(clk), .Q(fifo_array[879])
         );
  DFFPOSX1 fifo_array_reg_25__28_ ( .D(n2241), .CLK(clk), .Q(fifo_array[878])
         );
  DFFPOSX1 fifo_array_reg_25__27_ ( .D(n2240), .CLK(clk), .Q(fifo_array[877])
         );
  DFFPOSX1 fifo_array_reg_25__26_ ( .D(n2239), .CLK(clk), .Q(fifo_array[876])
         );
  DFFPOSX1 fifo_array_reg_25__25_ ( .D(n2238), .CLK(clk), .Q(fifo_array[875])
         );
  DFFPOSX1 fifo_array_reg_25__24_ ( .D(n2237), .CLK(clk), .Q(fifo_array[874])
         );
  DFFPOSX1 fifo_array_reg_25__23_ ( .D(n2236), .CLK(clk), .Q(fifo_array[873])
         );
  DFFPOSX1 fifo_array_reg_25__22_ ( .D(n2235), .CLK(clk), .Q(fifo_array[872])
         );
  DFFPOSX1 fifo_array_reg_25__21_ ( .D(n2234), .CLK(clk), .Q(fifo_array[871])
         );
  DFFPOSX1 fifo_array_reg_25__20_ ( .D(n2233), .CLK(clk), .Q(fifo_array[870])
         );
  DFFPOSX1 fifo_array_reg_25__19_ ( .D(n2232), .CLK(clk), .Q(fifo_array[869])
         );
  DFFPOSX1 fifo_array_reg_25__18_ ( .D(n2231), .CLK(clk), .Q(fifo_array[868])
         );
  DFFPOSX1 fifo_array_reg_25__17_ ( .D(n2230), .CLK(clk), .Q(fifo_array[867])
         );
  DFFPOSX1 fifo_array_reg_25__16_ ( .D(n2229), .CLK(clk), .Q(fifo_array[866])
         );
  DFFPOSX1 fifo_array_reg_25__15_ ( .D(n2228), .CLK(clk), .Q(fifo_array[865])
         );
  DFFPOSX1 fifo_array_reg_25__14_ ( .D(n2227), .CLK(clk), .Q(fifo_array[864])
         );
  DFFPOSX1 fifo_array_reg_25__13_ ( .D(n2226), .CLK(clk), .Q(fifo_array[863])
         );
  DFFPOSX1 fifo_array_reg_25__12_ ( .D(n2225), .CLK(clk), .Q(fifo_array[862])
         );
  DFFPOSX1 fifo_array_reg_25__11_ ( .D(n2224), .CLK(clk), .Q(fifo_array[861])
         );
  DFFPOSX1 fifo_array_reg_25__10_ ( .D(n2223), .CLK(clk), .Q(fifo_array[860])
         );
  DFFPOSX1 fifo_array_reg_25__9_ ( .D(n2222), .CLK(clk), .Q(fifo_array[859])
         );
  DFFPOSX1 fifo_array_reg_25__8_ ( .D(n2221), .CLK(clk), .Q(fifo_array[858])
         );
  DFFPOSX1 fifo_array_reg_25__7_ ( .D(n2220), .CLK(clk), .Q(fifo_array[857])
         );
  DFFPOSX1 fifo_array_reg_25__6_ ( .D(n2219), .CLK(clk), .Q(fifo_array[856])
         );
  DFFPOSX1 fifo_array_reg_25__5_ ( .D(n2218), .CLK(clk), .Q(fifo_array[855])
         );
  DFFPOSX1 fifo_array_reg_25__4_ ( .D(n2217), .CLK(clk), .Q(fifo_array[854])
         );
  DFFPOSX1 fifo_array_reg_25__3_ ( .D(n2216), .CLK(clk), .Q(fifo_array[853])
         );
  DFFPOSX1 fifo_array_reg_25__2_ ( .D(n2215), .CLK(clk), .Q(fifo_array[852])
         );
  DFFPOSX1 fifo_array_reg_25__1_ ( .D(n2214), .CLK(clk), .Q(fifo_array[851])
         );
  DFFPOSX1 fifo_array_reg_25__0_ ( .D(n2213), .CLK(clk), .Q(fifo_array[850])
         );
  DFFPOSX1 fifo_array_reg_24__33_ ( .D(n2212), .CLK(clk), .Q(fifo_array[849])
         );
  DFFPOSX1 fifo_array_reg_24__32_ ( .D(n2211), .CLK(clk), .Q(fifo_array[848])
         );
  DFFPOSX1 fifo_array_reg_24__31_ ( .D(n2210), .CLK(clk), .Q(fifo_array[847])
         );
  DFFPOSX1 fifo_array_reg_24__30_ ( .D(n2209), .CLK(clk), .Q(fifo_array[846])
         );
  DFFPOSX1 fifo_array_reg_24__29_ ( .D(n2208), .CLK(clk), .Q(fifo_array[845])
         );
  DFFPOSX1 fifo_array_reg_24__28_ ( .D(n2207), .CLK(clk), .Q(fifo_array[844])
         );
  DFFPOSX1 fifo_array_reg_24__27_ ( .D(n2206), .CLK(clk), .Q(fifo_array[843])
         );
  DFFPOSX1 fifo_array_reg_24__26_ ( .D(n2205), .CLK(clk), .Q(fifo_array[842])
         );
  DFFPOSX1 fifo_array_reg_24__25_ ( .D(n2204), .CLK(clk), .Q(fifo_array[841])
         );
  DFFPOSX1 fifo_array_reg_24__24_ ( .D(n2203), .CLK(clk), .Q(fifo_array[840])
         );
  DFFPOSX1 fifo_array_reg_24__23_ ( .D(n2202), .CLK(clk), .Q(fifo_array[839])
         );
  DFFPOSX1 fifo_array_reg_24__22_ ( .D(n2201), .CLK(clk), .Q(fifo_array[838])
         );
  DFFPOSX1 fifo_array_reg_24__21_ ( .D(n2200), .CLK(clk), .Q(fifo_array[837])
         );
  DFFPOSX1 fifo_array_reg_24__20_ ( .D(n2199), .CLK(clk), .Q(fifo_array[836])
         );
  DFFPOSX1 fifo_array_reg_24__19_ ( .D(n2198), .CLK(clk), .Q(fifo_array[835])
         );
  DFFPOSX1 fifo_array_reg_24__18_ ( .D(n2197), .CLK(clk), .Q(fifo_array[834])
         );
  DFFPOSX1 fifo_array_reg_24__17_ ( .D(n2196), .CLK(clk), .Q(fifo_array[833])
         );
  DFFPOSX1 fifo_array_reg_24__16_ ( .D(n2195), .CLK(clk), .Q(fifo_array[832])
         );
  DFFPOSX1 fifo_array_reg_24__15_ ( .D(n2194), .CLK(clk), .Q(fifo_array[831])
         );
  DFFPOSX1 fifo_array_reg_24__14_ ( .D(n2193), .CLK(clk), .Q(fifo_array[830])
         );
  DFFPOSX1 fifo_array_reg_24__13_ ( .D(n2192), .CLK(clk), .Q(fifo_array[829])
         );
  DFFPOSX1 fifo_array_reg_24__12_ ( .D(n2191), .CLK(clk), .Q(fifo_array[828])
         );
  DFFPOSX1 fifo_array_reg_24__11_ ( .D(n2190), .CLK(clk), .Q(fifo_array[827])
         );
  DFFPOSX1 fifo_array_reg_24__10_ ( .D(n2189), .CLK(clk), .Q(fifo_array[826])
         );
  DFFPOSX1 fifo_array_reg_24__9_ ( .D(n2188), .CLK(clk), .Q(fifo_array[825])
         );
  DFFPOSX1 fifo_array_reg_24__8_ ( .D(n2187), .CLK(clk), .Q(fifo_array[824])
         );
  DFFPOSX1 fifo_array_reg_24__7_ ( .D(n2186), .CLK(clk), .Q(fifo_array[823])
         );
  DFFPOSX1 fifo_array_reg_24__6_ ( .D(n2185), .CLK(clk), .Q(fifo_array[822])
         );
  DFFPOSX1 fifo_array_reg_24__5_ ( .D(n2184), .CLK(clk), .Q(fifo_array[821])
         );
  DFFPOSX1 fifo_array_reg_24__4_ ( .D(n2183), .CLK(clk), .Q(fifo_array[820])
         );
  DFFPOSX1 fifo_array_reg_24__3_ ( .D(n2182), .CLK(clk), .Q(fifo_array[819])
         );
  DFFPOSX1 fifo_array_reg_24__2_ ( .D(n2181), .CLK(clk), .Q(fifo_array[818])
         );
  DFFPOSX1 fifo_array_reg_24__1_ ( .D(n2180), .CLK(clk), .Q(fifo_array[817])
         );
  DFFPOSX1 fifo_array_reg_24__0_ ( .D(n2179), .CLK(clk), .Q(fifo_array[816])
         );
  DFFPOSX1 fifo_array_reg_23__33_ ( .D(n2178), .CLK(clk), .Q(fifo_array[815])
         );
  DFFPOSX1 fifo_array_reg_23__32_ ( .D(n2177), .CLK(clk), .Q(fifo_array[814])
         );
  DFFPOSX1 fifo_array_reg_23__31_ ( .D(n2176), .CLK(clk), .Q(fifo_array[813])
         );
  DFFPOSX1 fifo_array_reg_23__30_ ( .D(n2175), .CLK(clk), .Q(fifo_array[812])
         );
  DFFPOSX1 fifo_array_reg_23__29_ ( .D(n2174), .CLK(clk), .Q(fifo_array[811])
         );
  DFFPOSX1 fifo_array_reg_23__28_ ( .D(n2173), .CLK(clk), .Q(fifo_array[810])
         );
  DFFPOSX1 fifo_array_reg_23__27_ ( .D(n2172), .CLK(clk), .Q(fifo_array[809])
         );
  DFFPOSX1 fifo_array_reg_23__26_ ( .D(n2171), .CLK(clk), .Q(fifo_array[808])
         );
  DFFPOSX1 fifo_array_reg_23__25_ ( .D(n2170), .CLK(clk), .Q(fifo_array[807])
         );
  DFFPOSX1 fifo_array_reg_23__24_ ( .D(n2169), .CLK(clk), .Q(fifo_array[806])
         );
  DFFPOSX1 fifo_array_reg_23__23_ ( .D(n2168), .CLK(clk), .Q(fifo_array[805])
         );
  DFFPOSX1 fifo_array_reg_23__22_ ( .D(n2167), .CLK(clk), .Q(fifo_array[804])
         );
  DFFPOSX1 fifo_array_reg_23__21_ ( .D(n2166), .CLK(clk), .Q(fifo_array[803])
         );
  DFFPOSX1 fifo_array_reg_23__20_ ( .D(n2165), .CLK(clk), .Q(fifo_array[802])
         );
  DFFPOSX1 fifo_array_reg_23__19_ ( .D(n2164), .CLK(clk), .Q(fifo_array[801])
         );
  DFFPOSX1 fifo_array_reg_23__18_ ( .D(n2163), .CLK(clk), .Q(fifo_array[800])
         );
  DFFPOSX1 fifo_array_reg_23__17_ ( .D(n2162), .CLK(clk), .Q(fifo_array[799])
         );
  DFFPOSX1 fifo_array_reg_23__16_ ( .D(n2161), .CLK(clk), .Q(fifo_array[798])
         );
  DFFPOSX1 fifo_array_reg_23__15_ ( .D(n2160), .CLK(clk), .Q(fifo_array[797])
         );
  DFFPOSX1 fifo_array_reg_23__14_ ( .D(n2159), .CLK(clk), .Q(fifo_array[796])
         );
  DFFPOSX1 fifo_array_reg_23__13_ ( .D(n2158), .CLK(clk), .Q(fifo_array[795])
         );
  DFFPOSX1 fifo_array_reg_23__12_ ( .D(n2157), .CLK(clk), .Q(fifo_array[794])
         );
  DFFPOSX1 fifo_array_reg_23__11_ ( .D(n2156), .CLK(clk), .Q(fifo_array[793])
         );
  DFFPOSX1 fifo_array_reg_23__10_ ( .D(n2155), .CLK(clk), .Q(fifo_array[792])
         );
  DFFPOSX1 fifo_array_reg_23__9_ ( .D(n2154), .CLK(clk), .Q(fifo_array[791])
         );
  DFFPOSX1 fifo_array_reg_23__8_ ( .D(n2153), .CLK(clk), .Q(fifo_array[790])
         );
  DFFPOSX1 fifo_array_reg_23__7_ ( .D(n2152), .CLK(clk), .Q(fifo_array[789])
         );
  DFFPOSX1 fifo_array_reg_23__6_ ( .D(n2151), .CLK(clk), .Q(fifo_array[788])
         );
  DFFPOSX1 fifo_array_reg_23__5_ ( .D(n2150), .CLK(clk), .Q(fifo_array[787])
         );
  DFFPOSX1 fifo_array_reg_23__4_ ( .D(n2149), .CLK(clk), .Q(fifo_array[786])
         );
  DFFPOSX1 fifo_array_reg_23__3_ ( .D(n2148), .CLK(clk), .Q(fifo_array[785])
         );
  DFFPOSX1 fifo_array_reg_23__2_ ( .D(n2147), .CLK(clk), .Q(fifo_array[784])
         );
  DFFPOSX1 fifo_array_reg_23__1_ ( .D(n2146), .CLK(clk), .Q(fifo_array[783])
         );
  DFFPOSX1 fifo_array_reg_23__0_ ( .D(n2145), .CLK(clk), .Q(fifo_array[782])
         );
  DFFPOSX1 fifo_array_reg_22__33_ ( .D(n2144), .CLK(clk), .Q(fifo_array[781])
         );
  DFFPOSX1 fifo_array_reg_22__32_ ( .D(n2143), .CLK(clk), .Q(fifo_array[780])
         );
  DFFPOSX1 fifo_array_reg_22__31_ ( .D(n2142), .CLK(clk), .Q(fifo_array[779])
         );
  DFFPOSX1 fifo_array_reg_22__30_ ( .D(n2141), .CLK(clk), .Q(fifo_array[778])
         );
  DFFPOSX1 fifo_array_reg_22__29_ ( .D(n2140), .CLK(clk), .Q(fifo_array[777])
         );
  DFFPOSX1 fifo_array_reg_22__28_ ( .D(n2139), .CLK(clk), .Q(fifo_array[776])
         );
  DFFPOSX1 fifo_array_reg_22__27_ ( .D(n2138), .CLK(clk), .Q(fifo_array[775])
         );
  DFFPOSX1 fifo_array_reg_22__26_ ( .D(n2137), .CLK(clk), .Q(fifo_array[774])
         );
  DFFPOSX1 fifo_array_reg_22__25_ ( .D(n2136), .CLK(clk), .Q(fifo_array[773])
         );
  DFFPOSX1 fifo_array_reg_22__24_ ( .D(n2135), .CLK(clk), .Q(fifo_array[772])
         );
  DFFPOSX1 fifo_array_reg_22__23_ ( .D(n2134), .CLK(clk), .Q(fifo_array[771])
         );
  DFFPOSX1 fifo_array_reg_22__22_ ( .D(n2133), .CLK(clk), .Q(fifo_array[770])
         );
  DFFPOSX1 fifo_array_reg_22__21_ ( .D(n2132), .CLK(clk), .Q(fifo_array[769])
         );
  DFFPOSX1 fifo_array_reg_22__20_ ( .D(n2131), .CLK(clk), .Q(fifo_array[768])
         );
  DFFPOSX1 fifo_array_reg_22__19_ ( .D(n2130), .CLK(clk), .Q(fifo_array[767])
         );
  DFFPOSX1 fifo_array_reg_22__18_ ( .D(n2129), .CLK(clk), .Q(fifo_array[766])
         );
  DFFPOSX1 fifo_array_reg_22__17_ ( .D(n2128), .CLK(clk), .Q(fifo_array[765])
         );
  DFFPOSX1 fifo_array_reg_22__16_ ( .D(n2127), .CLK(clk), .Q(fifo_array[764])
         );
  DFFPOSX1 fifo_array_reg_22__15_ ( .D(n2126), .CLK(clk), .Q(fifo_array[763])
         );
  DFFPOSX1 fifo_array_reg_22__14_ ( .D(n2125), .CLK(clk), .Q(fifo_array[762])
         );
  DFFPOSX1 fifo_array_reg_22__13_ ( .D(n2124), .CLK(clk), .Q(fifo_array[761])
         );
  DFFPOSX1 fifo_array_reg_22__12_ ( .D(n2123), .CLK(clk), .Q(fifo_array[760])
         );
  DFFPOSX1 fifo_array_reg_22__11_ ( .D(n2122), .CLK(clk), .Q(fifo_array[759])
         );
  DFFPOSX1 fifo_array_reg_22__10_ ( .D(n2121), .CLK(clk), .Q(fifo_array[758])
         );
  DFFPOSX1 fifo_array_reg_22__9_ ( .D(n2120), .CLK(clk), .Q(fifo_array[757])
         );
  DFFPOSX1 fifo_array_reg_22__8_ ( .D(n2119), .CLK(clk), .Q(fifo_array[756])
         );
  DFFPOSX1 fifo_array_reg_22__7_ ( .D(n2118), .CLK(clk), .Q(fifo_array[755])
         );
  DFFPOSX1 fifo_array_reg_22__6_ ( .D(n2117), .CLK(clk), .Q(fifo_array[754])
         );
  DFFPOSX1 fifo_array_reg_22__5_ ( .D(n2116), .CLK(clk), .Q(fifo_array[753])
         );
  DFFPOSX1 fifo_array_reg_22__4_ ( .D(n2115), .CLK(clk), .Q(fifo_array[752])
         );
  DFFPOSX1 fifo_array_reg_22__3_ ( .D(n2114), .CLK(clk), .Q(fifo_array[751])
         );
  DFFPOSX1 fifo_array_reg_22__2_ ( .D(n2113), .CLK(clk), .Q(fifo_array[750])
         );
  DFFPOSX1 fifo_array_reg_22__1_ ( .D(n2112), .CLK(clk), .Q(fifo_array[749])
         );
  DFFPOSX1 fifo_array_reg_22__0_ ( .D(n2111), .CLK(clk), .Q(fifo_array[748])
         );
  DFFPOSX1 fifo_array_reg_21__33_ ( .D(n2110), .CLK(clk), .Q(fifo_array[747])
         );
  DFFPOSX1 fifo_array_reg_21__32_ ( .D(n2109), .CLK(clk), .Q(fifo_array[746])
         );
  DFFPOSX1 fifo_array_reg_21__31_ ( .D(n2108), .CLK(clk), .Q(fifo_array[745])
         );
  DFFPOSX1 fifo_array_reg_21__30_ ( .D(n2107), .CLK(clk), .Q(fifo_array[744])
         );
  DFFPOSX1 fifo_array_reg_21__29_ ( .D(n2106), .CLK(clk), .Q(fifo_array[743])
         );
  DFFPOSX1 fifo_array_reg_21__28_ ( .D(n2105), .CLK(clk), .Q(fifo_array[742])
         );
  DFFPOSX1 fifo_array_reg_21__27_ ( .D(n2104), .CLK(clk), .Q(fifo_array[741])
         );
  DFFPOSX1 fifo_array_reg_21__26_ ( .D(n2103), .CLK(clk), .Q(fifo_array[740])
         );
  DFFPOSX1 fifo_array_reg_21__25_ ( .D(n2102), .CLK(clk), .Q(fifo_array[739])
         );
  DFFPOSX1 fifo_array_reg_21__24_ ( .D(n2101), .CLK(clk), .Q(fifo_array[738])
         );
  DFFPOSX1 fifo_array_reg_21__23_ ( .D(n2100), .CLK(clk), .Q(fifo_array[737])
         );
  DFFPOSX1 fifo_array_reg_21__22_ ( .D(n2099), .CLK(clk), .Q(fifo_array[736])
         );
  DFFPOSX1 fifo_array_reg_21__21_ ( .D(n2098), .CLK(clk), .Q(fifo_array[735])
         );
  DFFPOSX1 fifo_array_reg_21__20_ ( .D(n2097), .CLK(clk), .Q(fifo_array[734])
         );
  DFFPOSX1 fifo_array_reg_21__19_ ( .D(n2096), .CLK(clk), .Q(fifo_array[733])
         );
  DFFPOSX1 fifo_array_reg_21__18_ ( .D(n2095), .CLK(clk), .Q(fifo_array[732])
         );
  DFFPOSX1 fifo_array_reg_21__17_ ( .D(n2094), .CLK(clk), .Q(fifo_array[731])
         );
  DFFPOSX1 fifo_array_reg_21__16_ ( .D(n2093), .CLK(clk), .Q(fifo_array[730])
         );
  DFFPOSX1 fifo_array_reg_21__15_ ( .D(n2092), .CLK(clk), .Q(fifo_array[729])
         );
  DFFPOSX1 fifo_array_reg_21__14_ ( .D(n2091), .CLK(clk), .Q(fifo_array[728])
         );
  DFFPOSX1 fifo_array_reg_21__13_ ( .D(n2090), .CLK(clk), .Q(fifo_array[727])
         );
  DFFPOSX1 fifo_array_reg_21__12_ ( .D(n2089), .CLK(clk), .Q(fifo_array[726])
         );
  DFFPOSX1 fifo_array_reg_21__11_ ( .D(n2088), .CLK(clk), .Q(fifo_array[725])
         );
  DFFPOSX1 fifo_array_reg_21__10_ ( .D(n2087), .CLK(clk), .Q(fifo_array[724])
         );
  DFFPOSX1 fifo_array_reg_21__9_ ( .D(n2086), .CLK(clk), .Q(fifo_array[723])
         );
  DFFPOSX1 fifo_array_reg_21__8_ ( .D(n2085), .CLK(clk), .Q(fifo_array[722])
         );
  DFFPOSX1 fifo_array_reg_21__7_ ( .D(n2084), .CLK(clk), .Q(fifo_array[721])
         );
  DFFPOSX1 fifo_array_reg_21__6_ ( .D(n2083), .CLK(clk), .Q(fifo_array[720])
         );
  DFFPOSX1 fifo_array_reg_21__5_ ( .D(n2082), .CLK(clk), .Q(fifo_array[719])
         );
  DFFPOSX1 fifo_array_reg_21__4_ ( .D(n2081), .CLK(clk), .Q(fifo_array[718])
         );
  DFFPOSX1 fifo_array_reg_21__3_ ( .D(n2080), .CLK(clk), .Q(fifo_array[717])
         );
  DFFPOSX1 fifo_array_reg_21__2_ ( .D(n2079), .CLK(clk), .Q(fifo_array[716])
         );
  DFFPOSX1 fifo_array_reg_21__1_ ( .D(n2078), .CLK(clk), .Q(fifo_array[715])
         );
  DFFPOSX1 fifo_array_reg_21__0_ ( .D(n2077), .CLK(clk), .Q(fifo_array[714])
         );
  DFFPOSX1 fifo_array_reg_20__33_ ( .D(n2076), .CLK(clk), .Q(fifo_array[713])
         );
  DFFPOSX1 fifo_array_reg_20__32_ ( .D(n2075), .CLK(clk), .Q(fifo_array[712])
         );
  DFFPOSX1 fifo_array_reg_20__31_ ( .D(n2074), .CLK(clk), .Q(fifo_array[711])
         );
  DFFPOSX1 fifo_array_reg_20__30_ ( .D(n2073), .CLK(clk), .Q(fifo_array[710])
         );
  DFFPOSX1 fifo_array_reg_20__29_ ( .D(n2072), .CLK(clk), .Q(fifo_array[709])
         );
  DFFPOSX1 fifo_array_reg_20__28_ ( .D(n2071), .CLK(clk), .Q(fifo_array[708])
         );
  DFFPOSX1 fifo_array_reg_20__27_ ( .D(n2070), .CLK(clk), .Q(fifo_array[707])
         );
  DFFPOSX1 fifo_array_reg_20__26_ ( .D(n2069), .CLK(clk), .Q(fifo_array[706])
         );
  DFFPOSX1 fifo_array_reg_20__25_ ( .D(n2068), .CLK(clk), .Q(fifo_array[705])
         );
  DFFPOSX1 fifo_array_reg_20__24_ ( .D(n2067), .CLK(clk), .Q(fifo_array[704])
         );
  DFFPOSX1 fifo_array_reg_20__23_ ( .D(n2066), .CLK(clk), .Q(fifo_array[703])
         );
  DFFPOSX1 fifo_array_reg_20__22_ ( .D(n2065), .CLK(clk), .Q(fifo_array[702])
         );
  DFFPOSX1 fifo_array_reg_20__21_ ( .D(n2064), .CLK(clk), .Q(fifo_array[701])
         );
  DFFPOSX1 fifo_array_reg_20__20_ ( .D(n2063), .CLK(clk), .Q(fifo_array[700])
         );
  DFFPOSX1 fifo_array_reg_20__19_ ( .D(n2062), .CLK(clk), .Q(fifo_array[699])
         );
  DFFPOSX1 fifo_array_reg_20__18_ ( .D(n2061), .CLK(clk), .Q(fifo_array[698])
         );
  DFFPOSX1 fifo_array_reg_20__17_ ( .D(n2060), .CLK(clk), .Q(fifo_array[697])
         );
  DFFPOSX1 fifo_array_reg_20__16_ ( .D(n2059), .CLK(clk), .Q(fifo_array[696])
         );
  DFFPOSX1 fifo_array_reg_20__15_ ( .D(n2058), .CLK(clk), .Q(fifo_array[695])
         );
  DFFPOSX1 fifo_array_reg_20__14_ ( .D(n2057), .CLK(clk), .Q(fifo_array[694])
         );
  DFFPOSX1 fifo_array_reg_20__13_ ( .D(n2056), .CLK(clk), .Q(fifo_array[693])
         );
  DFFPOSX1 fifo_array_reg_20__12_ ( .D(n2055), .CLK(clk), .Q(fifo_array[692])
         );
  DFFPOSX1 fifo_array_reg_20__11_ ( .D(n2054), .CLK(clk), .Q(fifo_array[691])
         );
  DFFPOSX1 fifo_array_reg_20__10_ ( .D(n2053), .CLK(clk), .Q(fifo_array[690])
         );
  DFFPOSX1 fifo_array_reg_20__9_ ( .D(n2052), .CLK(clk), .Q(fifo_array[689])
         );
  DFFPOSX1 fifo_array_reg_20__8_ ( .D(n2051), .CLK(clk), .Q(fifo_array[688])
         );
  DFFPOSX1 fifo_array_reg_20__7_ ( .D(n2050), .CLK(clk), .Q(fifo_array[687])
         );
  DFFPOSX1 fifo_array_reg_20__6_ ( .D(n2049), .CLK(clk), .Q(fifo_array[686])
         );
  DFFPOSX1 fifo_array_reg_20__5_ ( .D(n2048), .CLK(clk), .Q(fifo_array[685])
         );
  DFFPOSX1 fifo_array_reg_20__4_ ( .D(n2047), .CLK(clk), .Q(fifo_array[684])
         );
  DFFPOSX1 fifo_array_reg_20__3_ ( .D(n2046), .CLK(clk), .Q(fifo_array[683])
         );
  DFFPOSX1 fifo_array_reg_20__2_ ( .D(n2045), .CLK(clk), .Q(fifo_array[682])
         );
  DFFPOSX1 fifo_array_reg_20__1_ ( .D(n2044), .CLK(clk), .Q(fifo_array[681])
         );
  DFFPOSX1 fifo_array_reg_20__0_ ( .D(n2043), .CLK(clk), .Q(fifo_array[680])
         );
  DFFPOSX1 fifo_array_reg_19__33_ ( .D(n2042), .CLK(clk), .Q(fifo_array[679])
         );
  DFFPOSX1 fifo_array_reg_19__32_ ( .D(n2041), .CLK(clk), .Q(fifo_array[678])
         );
  DFFPOSX1 fifo_array_reg_19__31_ ( .D(n2040), .CLK(clk), .Q(fifo_array[677])
         );
  DFFPOSX1 fifo_array_reg_19__30_ ( .D(n2039), .CLK(clk), .Q(fifo_array[676])
         );
  DFFPOSX1 fifo_array_reg_19__29_ ( .D(n2038), .CLK(clk), .Q(fifo_array[675])
         );
  DFFPOSX1 fifo_array_reg_19__28_ ( .D(n2037), .CLK(clk), .Q(fifo_array[674])
         );
  DFFPOSX1 fifo_array_reg_19__27_ ( .D(n2036), .CLK(clk), .Q(fifo_array[673])
         );
  DFFPOSX1 fifo_array_reg_19__26_ ( .D(n2035), .CLK(clk), .Q(fifo_array[672])
         );
  DFFPOSX1 fifo_array_reg_19__25_ ( .D(n2034), .CLK(clk), .Q(fifo_array[671])
         );
  DFFPOSX1 fifo_array_reg_19__24_ ( .D(n2033), .CLK(clk), .Q(fifo_array[670])
         );
  DFFPOSX1 fifo_array_reg_19__23_ ( .D(n2032), .CLK(clk), .Q(fifo_array[669])
         );
  DFFPOSX1 fifo_array_reg_19__22_ ( .D(n2031), .CLK(clk), .Q(fifo_array[668])
         );
  DFFPOSX1 fifo_array_reg_19__21_ ( .D(n2030), .CLK(clk), .Q(fifo_array[667])
         );
  DFFPOSX1 fifo_array_reg_19__20_ ( .D(n2029), .CLK(clk), .Q(fifo_array[666])
         );
  DFFPOSX1 fifo_array_reg_19__19_ ( .D(n2028), .CLK(clk), .Q(fifo_array[665])
         );
  DFFPOSX1 fifo_array_reg_19__18_ ( .D(n2027), .CLK(clk), .Q(fifo_array[664])
         );
  DFFPOSX1 fifo_array_reg_19__17_ ( .D(n2026), .CLK(clk), .Q(fifo_array[663])
         );
  DFFPOSX1 fifo_array_reg_19__16_ ( .D(n2025), .CLK(clk), .Q(fifo_array[662])
         );
  DFFPOSX1 fifo_array_reg_19__15_ ( .D(n2024), .CLK(clk), .Q(fifo_array[661])
         );
  DFFPOSX1 fifo_array_reg_19__14_ ( .D(n2023), .CLK(clk), .Q(fifo_array[660])
         );
  DFFPOSX1 fifo_array_reg_19__13_ ( .D(n2022), .CLK(clk), .Q(fifo_array[659])
         );
  DFFPOSX1 fifo_array_reg_19__12_ ( .D(n2021), .CLK(clk), .Q(fifo_array[658])
         );
  DFFPOSX1 fifo_array_reg_19__11_ ( .D(n2020), .CLK(clk), .Q(fifo_array[657])
         );
  DFFPOSX1 fifo_array_reg_19__10_ ( .D(n2019), .CLK(clk), .Q(fifo_array[656])
         );
  DFFPOSX1 fifo_array_reg_19__9_ ( .D(n2018), .CLK(clk), .Q(fifo_array[655])
         );
  DFFPOSX1 fifo_array_reg_19__8_ ( .D(n2017), .CLK(clk), .Q(fifo_array[654])
         );
  DFFPOSX1 fifo_array_reg_19__7_ ( .D(n2016), .CLK(clk), .Q(fifo_array[653])
         );
  DFFPOSX1 fifo_array_reg_19__6_ ( .D(n2015), .CLK(clk), .Q(fifo_array[652])
         );
  DFFPOSX1 fifo_array_reg_19__5_ ( .D(n2014), .CLK(clk), .Q(fifo_array[651])
         );
  DFFPOSX1 fifo_array_reg_19__4_ ( .D(n2013), .CLK(clk), .Q(fifo_array[650])
         );
  DFFPOSX1 fifo_array_reg_19__3_ ( .D(n2012), .CLK(clk), .Q(fifo_array[649])
         );
  DFFPOSX1 fifo_array_reg_19__2_ ( .D(n2011), .CLK(clk), .Q(fifo_array[648])
         );
  DFFPOSX1 fifo_array_reg_19__1_ ( .D(n2010), .CLK(clk), .Q(fifo_array[647])
         );
  DFFPOSX1 fifo_array_reg_19__0_ ( .D(n2009), .CLK(clk), .Q(fifo_array[646])
         );
  DFFPOSX1 fifo_array_reg_18__33_ ( .D(n2008), .CLK(clk), .Q(fifo_array[645])
         );
  DFFPOSX1 fifo_array_reg_18__32_ ( .D(n2007), .CLK(clk), .Q(fifo_array[644])
         );
  DFFPOSX1 fifo_array_reg_18__31_ ( .D(n2006), .CLK(clk), .Q(fifo_array[643])
         );
  DFFPOSX1 fifo_array_reg_18__30_ ( .D(n2005), .CLK(clk), .Q(fifo_array[642])
         );
  DFFPOSX1 fifo_array_reg_18__29_ ( .D(n2004), .CLK(clk), .Q(fifo_array[641])
         );
  DFFPOSX1 fifo_array_reg_18__28_ ( .D(n2003), .CLK(clk), .Q(fifo_array[640])
         );
  DFFPOSX1 fifo_array_reg_18__27_ ( .D(n2002), .CLK(clk), .Q(fifo_array[639])
         );
  DFFPOSX1 fifo_array_reg_18__26_ ( .D(n2001), .CLK(clk), .Q(fifo_array[638])
         );
  DFFPOSX1 fifo_array_reg_18__25_ ( .D(n2000), .CLK(clk), .Q(fifo_array[637])
         );
  DFFPOSX1 fifo_array_reg_18__24_ ( .D(n1999), .CLK(clk), .Q(fifo_array[636])
         );
  DFFPOSX1 fifo_array_reg_18__23_ ( .D(n1998), .CLK(clk), .Q(fifo_array[635])
         );
  DFFPOSX1 fifo_array_reg_18__22_ ( .D(n1997), .CLK(clk), .Q(fifo_array[634])
         );
  DFFPOSX1 fifo_array_reg_18__21_ ( .D(n1996), .CLK(clk), .Q(fifo_array[633])
         );
  DFFPOSX1 fifo_array_reg_18__20_ ( .D(n1995), .CLK(clk), .Q(fifo_array[632])
         );
  DFFPOSX1 fifo_array_reg_18__19_ ( .D(n1994), .CLK(clk), .Q(fifo_array[631])
         );
  DFFPOSX1 fifo_array_reg_18__18_ ( .D(n1993), .CLK(clk), .Q(fifo_array[630])
         );
  DFFPOSX1 fifo_array_reg_18__17_ ( .D(n1992), .CLK(clk), .Q(fifo_array[629])
         );
  DFFPOSX1 fifo_array_reg_18__16_ ( .D(n1991), .CLK(clk), .Q(fifo_array[628])
         );
  DFFPOSX1 fifo_array_reg_18__15_ ( .D(n1990), .CLK(clk), .Q(fifo_array[627])
         );
  DFFPOSX1 fifo_array_reg_18__14_ ( .D(n1989), .CLK(clk), .Q(fifo_array[626])
         );
  DFFPOSX1 fifo_array_reg_18__13_ ( .D(n1988), .CLK(clk), .Q(fifo_array[625])
         );
  DFFPOSX1 fifo_array_reg_18__12_ ( .D(n1987), .CLK(clk), .Q(fifo_array[624])
         );
  DFFPOSX1 fifo_array_reg_18__11_ ( .D(n1986), .CLK(clk), .Q(fifo_array[623])
         );
  DFFPOSX1 fifo_array_reg_18__10_ ( .D(n1985), .CLK(clk), .Q(fifo_array[622])
         );
  DFFPOSX1 fifo_array_reg_18__9_ ( .D(n1984), .CLK(clk), .Q(fifo_array[621])
         );
  DFFPOSX1 fifo_array_reg_18__8_ ( .D(n1983), .CLK(clk), .Q(fifo_array[620])
         );
  DFFPOSX1 fifo_array_reg_18__7_ ( .D(n1982), .CLK(clk), .Q(fifo_array[619])
         );
  DFFPOSX1 fifo_array_reg_18__6_ ( .D(n1981), .CLK(clk), .Q(fifo_array[618])
         );
  DFFPOSX1 fifo_array_reg_18__5_ ( .D(n1980), .CLK(clk), .Q(fifo_array[617])
         );
  DFFPOSX1 fifo_array_reg_18__4_ ( .D(n1979), .CLK(clk), .Q(fifo_array[616])
         );
  DFFPOSX1 fifo_array_reg_18__3_ ( .D(n1978), .CLK(clk), .Q(fifo_array[615])
         );
  DFFPOSX1 fifo_array_reg_18__2_ ( .D(n1977), .CLK(clk), .Q(fifo_array[614])
         );
  DFFPOSX1 fifo_array_reg_18__1_ ( .D(n1976), .CLK(clk), .Q(fifo_array[613])
         );
  DFFPOSX1 fifo_array_reg_18__0_ ( .D(n1975), .CLK(clk), .Q(fifo_array[612])
         );
  DFFPOSX1 fifo_array_reg_17__33_ ( .D(n1974), .CLK(clk), .Q(fifo_array[611])
         );
  DFFPOSX1 fifo_array_reg_17__32_ ( .D(n1973), .CLK(clk), .Q(fifo_array[610])
         );
  DFFPOSX1 fifo_array_reg_17__31_ ( .D(n1972), .CLK(clk), .Q(fifo_array[609])
         );
  DFFPOSX1 fifo_array_reg_17__30_ ( .D(n1971), .CLK(clk), .Q(fifo_array[608])
         );
  DFFPOSX1 fifo_array_reg_17__29_ ( .D(n1970), .CLK(clk), .Q(fifo_array[607])
         );
  DFFPOSX1 fifo_array_reg_17__28_ ( .D(n1969), .CLK(clk), .Q(fifo_array[606])
         );
  DFFPOSX1 fifo_array_reg_17__27_ ( .D(n1968), .CLK(clk), .Q(fifo_array[605])
         );
  DFFPOSX1 fifo_array_reg_17__26_ ( .D(n1967), .CLK(clk), .Q(fifo_array[604])
         );
  DFFPOSX1 fifo_array_reg_17__25_ ( .D(n1966), .CLK(clk), .Q(fifo_array[603])
         );
  DFFPOSX1 fifo_array_reg_17__24_ ( .D(n1965), .CLK(clk), .Q(fifo_array[602])
         );
  DFFPOSX1 fifo_array_reg_17__23_ ( .D(n1964), .CLK(clk), .Q(fifo_array[601])
         );
  DFFPOSX1 fifo_array_reg_17__22_ ( .D(n1963), .CLK(clk), .Q(fifo_array[600])
         );
  DFFPOSX1 fifo_array_reg_17__21_ ( .D(n1962), .CLK(clk), .Q(fifo_array[599])
         );
  DFFPOSX1 fifo_array_reg_17__20_ ( .D(n1961), .CLK(clk), .Q(fifo_array[598])
         );
  DFFPOSX1 fifo_array_reg_17__19_ ( .D(n1960), .CLK(clk), .Q(fifo_array[597])
         );
  DFFPOSX1 fifo_array_reg_17__18_ ( .D(n1959), .CLK(clk), .Q(fifo_array[596])
         );
  DFFPOSX1 fifo_array_reg_17__17_ ( .D(n1958), .CLK(clk), .Q(fifo_array[595])
         );
  DFFPOSX1 fifo_array_reg_17__16_ ( .D(n1957), .CLK(clk), .Q(fifo_array[594])
         );
  DFFPOSX1 fifo_array_reg_17__15_ ( .D(n1956), .CLK(clk), .Q(fifo_array[593])
         );
  DFFPOSX1 fifo_array_reg_17__14_ ( .D(n1955), .CLK(clk), .Q(fifo_array[592])
         );
  DFFPOSX1 fifo_array_reg_17__13_ ( .D(n1954), .CLK(clk), .Q(fifo_array[591])
         );
  DFFPOSX1 fifo_array_reg_17__12_ ( .D(n1953), .CLK(clk), .Q(fifo_array[590])
         );
  DFFPOSX1 fifo_array_reg_17__11_ ( .D(n1952), .CLK(clk), .Q(fifo_array[589])
         );
  DFFPOSX1 fifo_array_reg_17__10_ ( .D(n1951), .CLK(clk), .Q(fifo_array[588])
         );
  DFFPOSX1 fifo_array_reg_17__9_ ( .D(n1950), .CLK(clk), .Q(fifo_array[587])
         );
  DFFPOSX1 fifo_array_reg_17__8_ ( .D(n1949), .CLK(clk), .Q(fifo_array[586])
         );
  DFFPOSX1 fifo_array_reg_17__7_ ( .D(n1948), .CLK(clk), .Q(fifo_array[585])
         );
  DFFPOSX1 fifo_array_reg_17__6_ ( .D(n1947), .CLK(clk), .Q(fifo_array[584])
         );
  DFFPOSX1 fifo_array_reg_17__5_ ( .D(n1946), .CLK(clk), .Q(fifo_array[583])
         );
  DFFPOSX1 fifo_array_reg_17__4_ ( .D(n1945), .CLK(clk), .Q(fifo_array[582])
         );
  DFFPOSX1 fifo_array_reg_17__3_ ( .D(n1944), .CLK(clk), .Q(fifo_array[581])
         );
  DFFPOSX1 fifo_array_reg_17__2_ ( .D(n1943), .CLK(clk), .Q(fifo_array[580])
         );
  DFFPOSX1 fifo_array_reg_17__1_ ( .D(n1942), .CLK(clk), .Q(fifo_array[579])
         );
  DFFPOSX1 fifo_array_reg_17__0_ ( .D(n1941), .CLK(clk), .Q(fifo_array[578])
         );
  DFFPOSX1 fifo_array_reg_16__33_ ( .D(n1940), .CLK(clk), .Q(fifo_array[577])
         );
  DFFPOSX1 fifo_array_reg_16__32_ ( .D(n1939), .CLK(clk), .Q(fifo_array[576])
         );
  DFFPOSX1 fifo_array_reg_16__31_ ( .D(n1938), .CLK(clk), .Q(fifo_array[575])
         );
  DFFPOSX1 fifo_array_reg_16__30_ ( .D(n1937), .CLK(clk), .Q(fifo_array[574])
         );
  DFFPOSX1 fifo_array_reg_16__29_ ( .D(n1936), .CLK(clk), .Q(fifo_array[573])
         );
  DFFPOSX1 fifo_array_reg_16__28_ ( .D(n1935), .CLK(clk), .Q(fifo_array[572])
         );
  DFFPOSX1 fifo_array_reg_16__27_ ( .D(n1934), .CLK(clk), .Q(fifo_array[571])
         );
  DFFPOSX1 fifo_array_reg_16__26_ ( .D(n1933), .CLK(clk), .Q(fifo_array[570])
         );
  DFFPOSX1 fifo_array_reg_16__25_ ( .D(n1932), .CLK(clk), .Q(fifo_array[569])
         );
  DFFPOSX1 fifo_array_reg_16__24_ ( .D(n1931), .CLK(clk), .Q(fifo_array[568])
         );
  DFFPOSX1 fifo_array_reg_16__23_ ( .D(n1930), .CLK(clk), .Q(fifo_array[567])
         );
  DFFPOSX1 fifo_array_reg_16__22_ ( .D(n1929), .CLK(clk), .Q(fifo_array[566])
         );
  DFFPOSX1 fifo_array_reg_16__21_ ( .D(n1928), .CLK(clk), .Q(fifo_array[565])
         );
  DFFPOSX1 fifo_array_reg_16__20_ ( .D(n1927), .CLK(clk), .Q(fifo_array[564])
         );
  DFFPOSX1 fifo_array_reg_16__19_ ( .D(n1926), .CLK(clk), .Q(fifo_array[563])
         );
  DFFPOSX1 fifo_array_reg_16__18_ ( .D(n1925), .CLK(clk), .Q(fifo_array[562])
         );
  DFFPOSX1 fifo_array_reg_16__17_ ( .D(n1924), .CLK(clk), .Q(fifo_array[561])
         );
  DFFPOSX1 fifo_array_reg_16__16_ ( .D(n1923), .CLK(clk), .Q(fifo_array[560])
         );
  DFFPOSX1 fifo_array_reg_16__15_ ( .D(n1922), .CLK(clk), .Q(fifo_array[559])
         );
  DFFPOSX1 fifo_array_reg_16__14_ ( .D(n1921), .CLK(clk), .Q(fifo_array[558])
         );
  DFFPOSX1 fifo_array_reg_16__13_ ( .D(n1920), .CLK(clk), .Q(fifo_array[557])
         );
  DFFPOSX1 fifo_array_reg_16__12_ ( .D(n1919), .CLK(clk), .Q(fifo_array[556])
         );
  DFFPOSX1 fifo_array_reg_16__11_ ( .D(n1918), .CLK(clk), .Q(fifo_array[555])
         );
  DFFPOSX1 fifo_array_reg_16__10_ ( .D(n1917), .CLK(clk), .Q(fifo_array[554])
         );
  DFFPOSX1 fifo_array_reg_16__9_ ( .D(n1916), .CLK(clk), .Q(fifo_array[553])
         );
  DFFPOSX1 fifo_array_reg_16__8_ ( .D(n1915), .CLK(clk), .Q(fifo_array[552])
         );
  DFFPOSX1 fifo_array_reg_16__7_ ( .D(n1914), .CLK(clk), .Q(fifo_array[551])
         );
  DFFPOSX1 fifo_array_reg_16__6_ ( .D(n1913), .CLK(clk), .Q(fifo_array[550])
         );
  DFFPOSX1 fifo_array_reg_16__5_ ( .D(n1912), .CLK(clk), .Q(fifo_array[549])
         );
  DFFPOSX1 fifo_array_reg_16__4_ ( .D(n1911), .CLK(clk), .Q(fifo_array[548])
         );
  DFFPOSX1 fifo_array_reg_16__3_ ( .D(n1910), .CLK(clk), .Q(fifo_array[547])
         );
  DFFPOSX1 fifo_array_reg_16__2_ ( .D(n1909), .CLK(clk), .Q(fifo_array[546])
         );
  DFFPOSX1 fifo_array_reg_16__1_ ( .D(n1908), .CLK(clk), .Q(fifo_array[545])
         );
  DFFPOSX1 fifo_array_reg_16__0_ ( .D(n1907), .CLK(clk), .Q(fifo_array[544])
         );
  DFFPOSX1 fifo_array_reg_15__33_ ( .D(n1906), .CLK(clk), .Q(fifo_array[543])
         );
  DFFPOSX1 fifo_array_reg_15__32_ ( .D(n1905), .CLK(clk), .Q(fifo_array[542])
         );
  DFFPOSX1 fifo_array_reg_15__31_ ( .D(n1904), .CLK(clk), .Q(fifo_array[541])
         );
  DFFPOSX1 fifo_array_reg_15__30_ ( .D(n1903), .CLK(clk), .Q(fifo_array[540])
         );
  DFFPOSX1 fifo_array_reg_15__29_ ( .D(n1902), .CLK(clk), .Q(fifo_array[539])
         );
  DFFPOSX1 fifo_array_reg_15__28_ ( .D(n1901), .CLK(clk), .Q(fifo_array[538])
         );
  DFFPOSX1 fifo_array_reg_15__27_ ( .D(n1900), .CLK(clk), .Q(fifo_array[537])
         );
  DFFPOSX1 fifo_array_reg_15__26_ ( .D(n1899), .CLK(clk), .Q(fifo_array[536])
         );
  DFFPOSX1 fifo_array_reg_15__25_ ( .D(n1898), .CLK(clk), .Q(fifo_array[535])
         );
  DFFPOSX1 fifo_array_reg_15__24_ ( .D(n1897), .CLK(clk), .Q(fifo_array[534])
         );
  DFFPOSX1 fifo_array_reg_15__23_ ( .D(n1896), .CLK(clk), .Q(fifo_array[533])
         );
  DFFPOSX1 fifo_array_reg_15__22_ ( .D(n1895), .CLK(clk), .Q(fifo_array[532])
         );
  DFFPOSX1 fifo_array_reg_15__21_ ( .D(n1894), .CLK(clk), .Q(fifo_array[531])
         );
  DFFPOSX1 fifo_array_reg_15__20_ ( .D(n1893), .CLK(clk), .Q(fifo_array[530])
         );
  DFFPOSX1 fifo_array_reg_15__19_ ( .D(n1892), .CLK(clk), .Q(fifo_array[529])
         );
  DFFPOSX1 fifo_array_reg_15__18_ ( .D(n1891), .CLK(clk), .Q(fifo_array[528])
         );
  DFFPOSX1 fifo_array_reg_15__17_ ( .D(n1890), .CLK(clk), .Q(fifo_array[527])
         );
  DFFPOSX1 fifo_array_reg_15__16_ ( .D(n1889), .CLK(clk), .Q(fifo_array[526])
         );
  DFFPOSX1 fifo_array_reg_15__15_ ( .D(n1888), .CLK(clk), .Q(fifo_array[525])
         );
  DFFPOSX1 fifo_array_reg_15__14_ ( .D(n1887), .CLK(clk), .Q(fifo_array[524])
         );
  DFFPOSX1 fifo_array_reg_15__13_ ( .D(n1886), .CLK(clk), .Q(fifo_array[523])
         );
  DFFPOSX1 fifo_array_reg_15__12_ ( .D(n1885), .CLK(clk), .Q(fifo_array[522])
         );
  DFFPOSX1 fifo_array_reg_15__11_ ( .D(n1884), .CLK(clk), .Q(fifo_array[521])
         );
  DFFPOSX1 fifo_array_reg_15__10_ ( .D(n1883), .CLK(clk), .Q(fifo_array[520])
         );
  DFFPOSX1 fifo_array_reg_15__9_ ( .D(n1882), .CLK(clk), .Q(fifo_array[519])
         );
  DFFPOSX1 fifo_array_reg_15__8_ ( .D(n1881), .CLK(clk), .Q(fifo_array[518])
         );
  DFFPOSX1 fifo_array_reg_15__7_ ( .D(n1880), .CLK(clk), .Q(fifo_array[517])
         );
  DFFPOSX1 fifo_array_reg_15__6_ ( .D(n1879), .CLK(clk), .Q(fifo_array[516])
         );
  DFFPOSX1 fifo_array_reg_15__5_ ( .D(n1878), .CLK(clk), .Q(fifo_array[515])
         );
  DFFPOSX1 fifo_array_reg_15__4_ ( .D(n1877), .CLK(clk), .Q(fifo_array[514])
         );
  DFFPOSX1 fifo_array_reg_15__3_ ( .D(n1876), .CLK(clk), .Q(fifo_array[513])
         );
  DFFPOSX1 fifo_array_reg_15__2_ ( .D(n1875), .CLK(clk), .Q(fifo_array[512])
         );
  DFFPOSX1 fifo_array_reg_15__1_ ( .D(n1874), .CLK(clk), .Q(fifo_array[511])
         );
  DFFPOSX1 fifo_array_reg_15__0_ ( .D(n1873), .CLK(clk), .Q(fifo_array[510])
         );
  DFFPOSX1 fifo_array_reg_14__33_ ( .D(n1872), .CLK(clk), .Q(fifo_array[509])
         );
  DFFPOSX1 fifo_array_reg_14__32_ ( .D(n1871), .CLK(clk), .Q(fifo_array[508])
         );
  DFFPOSX1 fifo_array_reg_14__31_ ( .D(n1870), .CLK(clk), .Q(fifo_array[507])
         );
  DFFPOSX1 fifo_array_reg_14__30_ ( .D(n1869), .CLK(clk), .Q(fifo_array[506])
         );
  DFFPOSX1 fifo_array_reg_14__29_ ( .D(n1868), .CLK(clk), .Q(fifo_array[505])
         );
  DFFPOSX1 fifo_array_reg_14__28_ ( .D(n1867), .CLK(clk), .Q(fifo_array[504])
         );
  DFFPOSX1 fifo_array_reg_14__27_ ( .D(n1866), .CLK(clk), .Q(fifo_array[503])
         );
  DFFPOSX1 fifo_array_reg_14__26_ ( .D(n1865), .CLK(clk), .Q(fifo_array[502])
         );
  DFFPOSX1 fifo_array_reg_14__25_ ( .D(n1864), .CLK(clk), .Q(fifo_array[501])
         );
  DFFPOSX1 fifo_array_reg_14__24_ ( .D(n1863), .CLK(clk), .Q(fifo_array[500])
         );
  DFFPOSX1 fifo_array_reg_14__23_ ( .D(n1862), .CLK(clk), .Q(fifo_array[499])
         );
  DFFPOSX1 fifo_array_reg_14__22_ ( .D(n1861), .CLK(clk), .Q(fifo_array[498])
         );
  DFFPOSX1 fifo_array_reg_14__21_ ( .D(n1860), .CLK(clk), .Q(fifo_array[497])
         );
  DFFPOSX1 fifo_array_reg_14__20_ ( .D(n1859), .CLK(clk), .Q(fifo_array[496])
         );
  DFFPOSX1 fifo_array_reg_14__19_ ( .D(n1858), .CLK(clk), .Q(fifo_array[495])
         );
  DFFPOSX1 fifo_array_reg_14__18_ ( .D(n1857), .CLK(clk), .Q(fifo_array[494])
         );
  DFFPOSX1 fifo_array_reg_14__17_ ( .D(n1856), .CLK(clk), .Q(fifo_array[493])
         );
  DFFPOSX1 fifo_array_reg_14__16_ ( .D(n1855), .CLK(clk), .Q(fifo_array[492])
         );
  DFFPOSX1 fifo_array_reg_14__15_ ( .D(n1854), .CLK(clk), .Q(fifo_array[491])
         );
  DFFPOSX1 fifo_array_reg_14__14_ ( .D(n1853), .CLK(clk), .Q(fifo_array[490])
         );
  DFFPOSX1 fifo_array_reg_14__13_ ( .D(n1852), .CLK(clk), .Q(fifo_array[489])
         );
  DFFPOSX1 fifo_array_reg_14__12_ ( .D(n1851), .CLK(clk), .Q(fifo_array[488])
         );
  DFFPOSX1 fifo_array_reg_14__11_ ( .D(n1850), .CLK(clk), .Q(fifo_array[487])
         );
  DFFPOSX1 fifo_array_reg_14__10_ ( .D(n1849), .CLK(clk), .Q(fifo_array[486])
         );
  DFFPOSX1 fifo_array_reg_14__9_ ( .D(n1848), .CLK(clk), .Q(fifo_array[485])
         );
  DFFPOSX1 fifo_array_reg_14__8_ ( .D(n1847), .CLK(clk), .Q(fifo_array[484])
         );
  DFFPOSX1 fifo_array_reg_14__7_ ( .D(n1846), .CLK(clk), .Q(fifo_array[483])
         );
  DFFPOSX1 fifo_array_reg_14__6_ ( .D(n1845), .CLK(clk), .Q(fifo_array[482])
         );
  DFFPOSX1 fifo_array_reg_14__5_ ( .D(n1844), .CLK(clk), .Q(fifo_array[481])
         );
  DFFPOSX1 fifo_array_reg_14__4_ ( .D(n1843), .CLK(clk), .Q(fifo_array[480])
         );
  DFFPOSX1 fifo_array_reg_14__3_ ( .D(n1842), .CLK(clk), .Q(fifo_array[479])
         );
  DFFPOSX1 fifo_array_reg_14__2_ ( .D(n1841), .CLK(clk), .Q(fifo_array[478])
         );
  DFFPOSX1 fifo_array_reg_14__1_ ( .D(n1840), .CLK(clk), .Q(fifo_array[477])
         );
  DFFPOSX1 fifo_array_reg_14__0_ ( .D(n1839), .CLK(clk), .Q(fifo_array[476])
         );
  DFFPOSX1 fifo_array_reg_13__33_ ( .D(n1838), .CLK(clk), .Q(fifo_array[475])
         );
  DFFPOSX1 fifo_array_reg_13__32_ ( .D(n1837), .CLK(clk), .Q(fifo_array[474])
         );
  DFFPOSX1 fifo_array_reg_13__31_ ( .D(n1836), .CLK(clk), .Q(fifo_array[473])
         );
  DFFPOSX1 fifo_array_reg_13__30_ ( .D(n1835), .CLK(clk), .Q(fifo_array[472])
         );
  DFFPOSX1 fifo_array_reg_13__29_ ( .D(n1834), .CLK(clk), .Q(fifo_array[471])
         );
  DFFPOSX1 fifo_array_reg_13__28_ ( .D(n1833), .CLK(clk), .Q(fifo_array[470])
         );
  DFFPOSX1 fifo_array_reg_13__27_ ( .D(n1832), .CLK(clk), .Q(fifo_array[469])
         );
  DFFPOSX1 fifo_array_reg_13__26_ ( .D(n1831), .CLK(clk), .Q(fifo_array[468])
         );
  DFFPOSX1 fifo_array_reg_13__25_ ( .D(n1830), .CLK(clk), .Q(fifo_array[467])
         );
  DFFPOSX1 fifo_array_reg_13__24_ ( .D(n1829), .CLK(clk), .Q(fifo_array[466])
         );
  DFFPOSX1 fifo_array_reg_13__23_ ( .D(n1828), .CLK(clk), .Q(fifo_array[465])
         );
  DFFPOSX1 fifo_array_reg_13__22_ ( .D(n1827), .CLK(clk), .Q(fifo_array[464])
         );
  DFFPOSX1 fifo_array_reg_13__21_ ( .D(n1826), .CLK(clk), .Q(fifo_array[463])
         );
  DFFPOSX1 fifo_array_reg_13__20_ ( .D(n1825), .CLK(clk), .Q(fifo_array[462])
         );
  DFFPOSX1 fifo_array_reg_13__19_ ( .D(n1824), .CLK(clk), .Q(fifo_array[461])
         );
  DFFPOSX1 fifo_array_reg_13__18_ ( .D(n1823), .CLK(clk), .Q(fifo_array[460])
         );
  DFFPOSX1 fifo_array_reg_13__17_ ( .D(n1822), .CLK(clk), .Q(fifo_array[459])
         );
  DFFPOSX1 fifo_array_reg_13__16_ ( .D(n1821), .CLK(clk), .Q(fifo_array[458])
         );
  DFFPOSX1 fifo_array_reg_13__15_ ( .D(n1820), .CLK(clk), .Q(fifo_array[457])
         );
  DFFPOSX1 fifo_array_reg_13__14_ ( .D(n1819), .CLK(clk), .Q(fifo_array[456])
         );
  DFFPOSX1 fifo_array_reg_13__13_ ( .D(n1818), .CLK(clk), .Q(fifo_array[455])
         );
  DFFPOSX1 fifo_array_reg_13__12_ ( .D(n1817), .CLK(clk), .Q(fifo_array[454])
         );
  DFFPOSX1 fifo_array_reg_13__11_ ( .D(n1816), .CLK(clk), .Q(fifo_array[453])
         );
  DFFPOSX1 fifo_array_reg_13__10_ ( .D(n1815), .CLK(clk), .Q(fifo_array[452])
         );
  DFFPOSX1 fifo_array_reg_13__9_ ( .D(n1814), .CLK(clk), .Q(fifo_array[451])
         );
  DFFPOSX1 fifo_array_reg_13__8_ ( .D(n1813), .CLK(clk), .Q(fifo_array[450])
         );
  DFFPOSX1 fifo_array_reg_13__7_ ( .D(n1812), .CLK(clk), .Q(fifo_array[449])
         );
  DFFPOSX1 fifo_array_reg_13__6_ ( .D(n1811), .CLK(clk), .Q(fifo_array[448])
         );
  DFFPOSX1 fifo_array_reg_13__5_ ( .D(n1810), .CLK(clk), .Q(fifo_array[447])
         );
  DFFPOSX1 fifo_array_reg_13__4_ ( .D(n1809), .CLK(clk), .Q(fifo_array[446])
         );
  DFFPOSX1 fifo_array_reg_13__3_ ( .D(n1808), .CLK(clk), .Q(fifo_array[445])
         );
  DFFPOSX1 fifo_array_reg_13__2_ ( .D(n1807), .CLK(clk), .Q(fifo_array[444])
         );
  DFFPOSX1 fifo_array_reg_13__1_ ( .D(n1806), .CLK(clk), .Q(fifo_array[443])
         );
  DFFPOSX1 fifo_array_reg_13__0_ ( .D(n1805), .CLK(clk), .Q(fifo_array[442])
         );
  DFFPOSX1 fifo_array_reg_12__33_ ( .D(n1804), .CLK(clk), .Q(fifo_array[441])
         );
  DFFPOSX1 fifo_array_reg_12__32_ ( .D(n1803), .CLK(clk), .Q(fifo_array[440])
         );
  DFFPOSX1 fifo_array_reg_12__31_ ( .D(n1802), .CLK(clk), .Q(fifo_array[439])
         );
  DFFPOSX1 fifo_array_reg_12__30_ ( .D(n1801), .CLK(clk), .Q(fifo_array[438])
         );
  DFFPOSX1 fifo_array_reg_12__29_ ( .D(n1800), .CLK(clk), .Q(fifo_array[437])
         );
  DFFPOSX1 fifo_array_reg_12__28_ ( .D(n1799), .CLK(clk), .Q(fifo_array[436])
         );
  DFFPOSX1 fifo_array_reg_12__27_ ( .D(n1798), .CLK(clk), .Q(fifo_array[435])
         );
  DFFPOSX1 fifo_array_reg_12__26_ ( .D(n1797), .CLK(clk), .Q(fifo_array[434])
         );
  DFFPOSX1 fifo_array_reg_12__25_ ( .D(n1796), .CLK(clk), .Q(fifo_array[433])
         );
  DFFPOSX1 fifo_array_reg_12__24_ ( .D(n1795), .CLK(clk), .Q(fifo_array[432])
         );
  DFFPOSX1 fifo_array_reg_12__23_ ( .D(n1794), .CLK(clk), .Q(fifo_array[431])
         );
  DFFPOSX1 fifo_array_reg_12__22_ ( .D(n1793), .CLK(clk), .Q(fifo_array[430])
         );
  DFFPOSX1 fifo_array_reg_12__21_ ( .D(n1792), .CLK(clk), .Q(fifo_array[429])
         );
  DFFPOSX1 fifo_array_reg_12__20_ ( .D(n1791), .CLK(clk), .Q(fifo_array[428])
         );
  DFFPOSX1 fifo_array_reg_12__19_ ( .D(n1790), .CLK(clk), .Q(fifo_array[427])
         );
  DFFPOSX1 fifo_array_reg_12__18_ ( .D(n1789), .CLK(clk), .Q(fifo_array[426])
         );
  DFFPOSX1 fifo_array_reg_12__17_ ( .D(n1788), .CLK(clk), .Q(fifo_array[425])
         );
  DFFPOSX1 fifo_array_reg_12__16_ ( .D(n1787), .CLK(clk), .Q(fifo_array[424])
         );
  DFFPOSX1 fifo_array_reg_12__15_ ( .D(n1786), .CLK(clk), .Q(fifo_array[423])
         );
  DFFPOSX1 fifo_array_reg_12__14_ ( .D(n1785), .CLK(clk), .Q(fifo_array[422])
         );
  DFFPOSX1 fifo_array_reg_12__13_ ( .D(n1784), .CLK(clk), .Q(fifo_array[421])
         );
  DFFPOSX1 fifo_array_reg_12__12_ ( .D(n1783), .CLK(clk), .Q(fifo_array[420])
         );
  DFFPOSX1 fifo_array_reg_12__11_ ( .D(n1782), .CLK(clk), .Q(fifo_array[419])
         );
  DFFPOSX1 fifo_array_reg_12__10_ ( .D(n1781), .CLK(clk), .Q(fifo_array[418])
         );
  DFFPOSX1 fifo_array_reg_12__9_ ( .D(n1780), .CLK(clk), .Q(fifo_array[417])
         );
  DFFPOSX1 fifo_array_reg_12__8_ ( .D(n1779), .CLK(clk), .Q(fifo_array[416])
         );
  DFFPOSX1 fifo_array_reg_12__7_ ( .D(n1778), .CLK(clk), .Q(fifo_array[415])
         );
  DFFPOSX1 fifo_array_reg_12__6_ ( .D(n1777), .CLK(clk), .Q(fifo_array[414])
         );
  DFFPOSX1 fifo_array_reg_12__5_ ( .D(n1776), .CLK(clk), .Q(fifo_array[413])
         );
  DFFPOSX1 fifo_array_reg_12__4_ ( .D(n1775), .CLK(clk), .Q(fifo_array[412])
         );
  DFFPOSX1 fifo_array_reg_12__3_ ( .D(n1774), .CLK(clk), .Q(fifo_array[411])
         );
  DFFPOSX1 fifo_array_reg_12__2_ ( .D(n1773), .CLK(clk), .Q(fifo_array[410])
         );
  DFFPOSX1 fifo_array_reg_12__1_ ( .D(n1772), .CLK(clk), .Q(fifo_array[409])
         );
  DFFPOSX1 fifo_array_reg_12__0_ ( .D(n1771), .CLK(clk), .Q(fifo_array[408])
         );
  DFFPOSX1 fifo_array_reg_11__33_ ( .D(n1770), .CLK(clk), .Q(fifo_array[407])
         );
  DFFPOSX1 fifo_array_reg_11__32_ ( .D(n1769), .CLK(clk), .Q(fifo_array[406])
         );
  DFFPOSX1 fifo_array_reg_11__31_ ( .D(n1768), .CLK(clk), .Q(fifo_array[405])
         );
  DFFPOSX1 fifo_array_reg_11__30_ ( .D(n1767), .CLK(clk), .Q(fifo_array[404])
         );
  DFFPOSX1 fifo_array_reg_11__29_ ( .D(n1766), .CLK(clk), .Q(fifo_array[403])
         );
  DFFPOSX1 fifo_array_reg_11__28_ ( .D(n1765), .CLK(clk), .Q(fifo_array[402])
         );
  DFFPOSX1 fifo_array_reg_11__27_ ( .D(n1764), .CLK(clk), .Q(fifo_array[401])
         );
  DFFPOSX1 fifo_array_reg_11__26_ ( .D(n1763), .CLK(clk), .Q(fifo_array[400])
         );
  DFFPOSX1 fifo_array_reg_11__25_ ( .D(n1762), .CLK(clk), .Q(fifo_array[399])
         );
  DFFPOSX1 fifo_array_reg_11__24_ ( .D(n1761), .CLK(clk), .Q(fifo_array[398])
         );
  DFFPOSX1 fifo_array_reg_11__23_ ( .D(n1760), .CLK(clk), .Q(fifo_array[397])
         );
  DFFPOSX1 fifo_array_reg_11__22_ ( .D(n1759), .CLK(clk), .Q(fifo_array[396])
         );
  DFFPOSX1 fifo_array_reg_11__21_ ( .D(n1758), .CLK(clk), .Q(fifo_array[395])
         );
  DFFPOSX1 fifo_array_reg_11__20_ ( .D(n1757), .CLK(clk), .Q(fifo_array[394])
         );
  DFFPOSX1 fifo_array_reg_11__19_ ( .D(n1756), .CLK(clk), .Q(fifo_array[393])
         );
  DFFPOSX1 fifo_array_reg_11__18_ ( .D(n1755), .CLK(clk), .Q(fifo_array[392])
         );
  DFFPOSX1 fifo_array_reg_11__17_ ( .D(n1754), .CLK(clk), .Q(fifo_array[391])
         );
  DFFPOSX1 fifo_array_reg_11__16_ ( .D(n1753), .CLK(clk), .Q(fifo_array[390])
         );
  DFFPOSX1 fifo_array_reg_11__15_ ( .D(n1752), .CLK(clk), .Q(fifo_array[389])
         );
  DFFPOSX1 fifo_array_reg_11__14_ ( .D(n1751), .CLK(clk), .Q(fifo_array[388])
         );
  DFFPOSX1 fifo_array_reg_11__13_ ( .D(n1750), .CLK(clk), .Q(fifo_array[387])
         );
  DFFPOSX1 fifo_array_reg_11__12_ ( .D(n1749), .CLK(clk), .Q(fifo_array[386])
         );
  DFFPOSX1 fifo_array_reg_11__11_ ( .D(n1748), .CLK(clk), .Q(fifo_array[385])
         );
  DFFPOSX1 fifo_array_reg_11__10_ ( .D(n1747), .CLK(clk), .Q(fifo_array[384])
         );
  DFFPOSX1 fifo_array_reg_11__9_ ( .D(n1746), .CLK(clk), .Q(fifo_array[383])
         );
  DFFPOSX1 fifo_array_reg_11__8_ ( .D(n1745), .CLK(clk), .Q(fifo_array[382])
         );
  DFFPOSX1 fifo_array_reg_11__7_ ( .D(n1744), .CLK(clk), .Q(fifo_array[381])
         );
  DFFPOSX1 fifo_array_reg_11__6_ ( .D(n1743), .CLK(clk), .Q(fifo_array[380])
         );
  DFFPOSX1 fifo_array_reg_11__5_ ( .D(n1742), .CLK(clk), .Q(fifo_array[379])
         );
  DFFPOSX1 fifo_array_reg_11__4_ ( .D(n1741), .CLK(clk), .Q(fifo_array[378])
         );
  DFFPOSX1 fifo_array_reg_11__3_ ( .D(n1740), .CLK(clk), .Q(fifo_array[377])
         );
  DFFPOSX1 fifo_array_reg_11__2_ ( .D(n1739), .CLK(clk), .Q(fifo_array[376])
         );
  DFFPOSX1 fifo_array_reg_11__1_ ( .D(n1738), .CLK(clk), .Q(fifo_array[375])
         );
  DFFPOSX1 fifo_array_reg_11__0_ ( .D(n1737), .CLK(clk), .Q(fifo_array[374])
         );
  DFFPOSX1 fifo_array_reg_10__33_ ( .D(n1736), .CLK(clk), .Q(fifo_array[373])
         );
  DFFPOSX1 fifo_array_reg_10__32_ ( .D(n1735), .CLK(clk), .Q(fifo_array[372])
         );
  DFFPOSX1 fifo_array_reg_10__31_ ( .D(n1734), .CLK(clk), .Q(fifo_array[371])
         );
  DFFPOSX1 fifo_array_reg_10__30_ ( .D(n1733), .CLK(clk), .Q(fifo_array[370])
         );
  DFFPOSX1 fifo_array_reg_10__29_ ( .D(n1732), .CLK(clk), .Q(fifo_array[369])
         );
  DFFPOSX1 fifo_array_reg_10__28_ ( .D(n1731), .CLK(clk), .Q(fifo_array[368])
         );
  DFFPOSX1 fifo_array_reg_10__27_ ( .D(n1730), .CLK(clk), .Q(fifo_array[367])
         );
  DFFPOSX1 fifo_array_reg_10__26_ ( .D(n1729), .CLK(clk), .Q(fifo_array[366])
         );
  DFFPOSX1 fifo_array_reg_10__25_ ( .D(n1728), .CLK(clk), .Q(fifo_array[365])
         );
  DFFPOSX1 fifo_array_reg_10__24_ ( .D(n1727), .CLK(clk), .Q(fifo_array[364])
         );
  DFFPOSX1 fifo_array_reg_10__23_ ( .D(n1726), .CLK(clk), .Q(fifo_array[363])
         );
  DFFPOSX1 fifo_array_reg_10__22_ ( .D(n1725), .CLK(clk), .Q(fifo_array[362])
         );
  DFFPOSX1 fifo_array_reg_10__21_ ( .D(n1724), .CLK(clk), .Q(fifo_array[361])
         );
  DFFPOSX1 fifo_array_reg_10__20_ ( .D(n1723), .CLK(clk), .Q(fifo_array[360])
         );
  DFFPOSX1 fifo_array_reg_10__19_ ( .D(n1722), .CLK(clk), .Q(fifo_array[359])
         );
  DFFPOSX1 fifo_array_reg_10__18_ ( .D(n1721), .CLK(clk), .Q(fifo_array[358])
         );
  DFFPOSX1 fifo_array_reg_10__17_ ( .D(n1720), .CLK(clk), .Q(fifo_array[357])
         );
  DFFPOSX1 fifo_array_reg_10__16_ ( .D(n1719), .CLK(clk), .Q(fifo_array[356])
         );
  DFFPOSX1 fifo_array_reg_10__15_ ( .D(n1718), .CLK(clk), .Q(fifo_array[355])
         );
  DFFPOSX1 fifo_array_reg_10__14_ ( .D(n1717), .CLK(clk), .Q(fifo_array[354])
         );
  DFFPOSX1 fifo_array_reg_10__13_ ( .D(n1716), .CLK(clk), .Q(fifo_array[353])
         );
  DFFPOSX1 fifo_array_reg_10__12_ ( .D(n1715), .CLK(clk), .Q(fifo_array[352])
         );
  DFFPOSX1 fifo_array_reg_10__11_ ( .D(n1714), .CLK(clk), .Q(fifo_array[351])
         );
  DFFPOSX1 fifo_array_reg_10__10_ ( .D(n1713), .CLK(clk), .Q(fifo_array[350])
         );
  DFFPOSX1 fifo_array_reg_10__9_ ( .D(n1712), .CLK(clk), .Q(fifo_array[349])
         );
  DFFPOSX1 fifo_array_reg_10__8_ ( .D(n1711), .CLK(clk), .Q(fifo_array[348])
         );
  DFFPOSX1 fifo_array_reg_10__7_ ( .D(n1710), .CLK(clk), .Q(fifo_array[347])
         );
  DFFPOSX1 fifo_array_reg_10__6_ ( .D(n1709), .CLK(clk), .Q(fifo_array[346])
         );
  DFFPOSX1 fifo_array_reg_10__5_ ( .D(n1708), .CLK(clk), .Q(fifo_array[345])
         );
  DFFPOSX1 fifo_array_reg_10__4_ ( .D(n1707), .CLK(clk), .Q(fifo_array[344])
         );
  DFFPOSX1 fifo_array_reg_10__3_ ( .D(n1706), .CLK(clk), .Q(fifo_array[343])
         );
  DFFPOSX1 fifo_array_reg_10__2_ ( .D(n1705), .CLK(clk), .Q(fifo_array[342])
         );
  DFFPOSX1 fifo_array_reg_10__1_ ( .D(n1704), .CLK(clk), .Q(fifo_array[341])
         );
  DFFPOSX1 fifo_array_reg_10__0_ ( .D(n1703), .CLK(clk), .Q(fifo_array[340])
         );
  DFFPOSX1 fifo_array_reg_9__33_ ( .D(n1702), .CLK(clk), .Q(fifo_array[339])
         );
  DFFPOSX1 fifo_array_reg_9__32_ ( .D(n1701), .CLK(clk), .Q(fifo_array[338])
         );
  DFFPOSX1 fifo_array_reg_9__31_ ( .D(n1700), .CLK(clk), .Q(fifo_array[337])
         );
  DFFPOSX1 fifo_array_reg_9__30_ ( .D(n1699), .CLK(clk), .Q(fifo_array[336])
         );
  DFFPOSX1 fifo_array_reg_9__29_ ( .D(n1698), .CLK(clk), .Q(fifo_array[335])
         );
  DFFPOSX1 fifo_array_reg_9__28_ ( .D(n1697), .CLK(clk), .Q(fifo_array[334])
         );
  DFFPOSX1 fifo_array_reg_9__27_ ( .D(n1696), .CLK(clk), .Q(fifo_array[333])
         );
  DFFPOSX1 fifo_array_reg_9__26_ ( .D(n1695), .CLK(clk), .Q(fifo_array[332])
         );
  DFFPOSX1 fifo_array_reg_9__25_ ( .D(n1694), .CLK(clk), .Q(fifo_array[331])
         );
  DFFPOSX1 fifo_array_reg_9__24_ ( .D(n1693), .CLK(clk), .Q(fifo_array[330])
         );
  DFFPOSX1 fifo_array_reg_9__23_ ( .D(n1692), .CLK(clk), .Q(fifo_array[329])
         );
  DFFPOSX1 fifo_array_reg_9__22_ ( .D(n1691), .CLK(clk), .Q(fifo_array[328])
         );
  DFFPOSX1 fifo_array_reg_9__21_ ( .D(n1690), .CLK(clk), .Q(fifo_array[327])
         );
  DFFPOSX1 fifo_array_reg_9__20_ ( .D(n1689), .CLK(clk), .Q(fifo_array[326])
         );
  DFFPOSX1 fifo_array_reg_9__19_ ( .D(n1688), .CLK(clk), .Q(fifo_array[325])
         );
  DFFPOSX1 fifo_array_reg_9__18_ ( .D(n1687), .CLK(clk), .Q(fifo_array[324])
         );
  DFFPOSX1 fifo_array_reg_9__17_ ( .D(n1686), .CLK(clk), .Q(fifo_array[323])
         );
  DFFPOSX1 fifo_array_reg_9__16_ ( .D(n1685), .CLK(clk), .Q(fifo_array[322])
         );
  DFFPOSX1 fifo_array_reg_9__15_ ( .D(n1684), .CLK(clk), .Q(fifo_array[321])
         );
  DFFPOSX1 fifo_array_reg_9__14_ ( .D(n1683), .CLK(clk), .Q(fifo_array[320])
         );
  DFFPOSX1 fifo_array_reg_9__13_ ( .D(n1682), .CLK(clk), .Q(fifo_array[319])
         );
  DFFPOSX1 fifo_array_reg_9__12_ ( .D(n1681), .CLK(clk), .Q(fifo_array[318])
         );
  DFFPOSX1 fifo_array_reg_9__11_ ( .D(n1680), .CLK(clk), .Q(fifo_array[317])
         );
  DFFPOSX1 fifo_array_reg_9__10_ ( .D(n1679), .CLK(clk), .Q(fifo_array[316])
         );
  DFFPOSX1 fifo_array_reg_9__9_ ( .D(n1678), .CLK(clk), .Q(fifo_array[315]) );
  DFFPOSX1 fifo_array_reg_9__8_ ( .D(n1677), .CLK(clk), .Q(fifo_array[314]) );
  DFFPOSX1 fifo_array_reg_9__7_ ( .D(n1676), .CLK(clk), .Q(fifo_array[313]) );
  DFFPOSX1 fifo_array_reg_9__6_ ( .D(n1675), .CLK(clk), .Q(fifo_array[312]) );
  DFFPOSX1 fifo_array_reg_9__5_ ( .D(n1674), .CLK(clk), .Q(fifo_array[311]) );
  DFFPOSX1 fifo_array_reg_9__4_ ( .D(n1673), .CLK(clk), .Q(fifo_array[310]) );
  DFFPOSX1 fifo_array_reg_9__3_ ( .D(n1672), .CLK(clk), .Q(fifo_array[309]) );
  DFFPOSX1 fifo_array_reg_9__2_ ( .D(n1671), .CLK(clk), .Q(fifo_array[308]) );
  DFFPOSX1 fifo_array_reg_9__1_ ( .D(n1670), .CLK(clk), .Q(fifo_array[307]) );
  DFFPOSX1 fifo_array_reg_9__0_ ( .D(n1669), .CLK(clk), .Q(fifo_array[306]) );
  DFFPOSX1 fifo_array_reg_8__33_ ( .D(n1668), .CLK(clk), .Q(fifo_array[305])
         );
  DFFPOSX1 fifo_array_reg_8__32_ ( .D(n1667), .CLK(clk), .Q(fifo_array[304])
         );
  DFFPOSX1 fifo_array_reg_8__31_ ( .D(n1666), .CLK(clk), .Q(fifo_array[303])
         );
  DFFPOSX1 fifo_array_reg_8__30_ ( .D(n1665), .CLK(clk), .Q(fifo_array[302])
         );
  DFFPOSX1 fifo_array_reg_8__29_ ( .D(n1664), .CLK(clk), .Q(fifo_array[301])
         );
  DFFPOSX1 fifo_array_reg_8__28_ ( .D(n1663), .CLK(clk), .Q(fifo_array[300])
         );
  DFFPOSX1 fifo_array_reg_8__27_ ( .D(n1662), .CLK(clk), .Q(fifo_array[299])
         );
  DFFPOSX1 fifo_array_reg_8__26_ ( .D(n1661), .CLK(clk), .Q(fifo_array[298])
         );
  DFFPOSX1 fifo_array_reg_8__25_ ( .D(n1660), .CLK(clk), .Q(fifo_array[297])
         );
  DFFPOSX1 fifo_array_reg_8__24_ ( .D(n1659), .CLK(clk), .Q(fifo_array[296])
         );
  DFFPOSX1 fifo_array_reg_8__23_ ( .D(n1658), .CLK(clk), .Q(fifo_array[295])
         );
  DFFPOSX1 fifo_array_reg_8__22_ ( .D(n1657), .CLK(clk), .Q(fifo_array[294])
         );
  DFFPOSX1 fifo_array_reg_8__21_ ( .D(n1656), .CLK(clk), .Q(fifo_array[293])
         );
  DFFPOSX1 fifo_array_reg_8__20_ ( .D(n1655), .CLK(clk), .Q(fifo_array[292])
         );
  DFFPOSX1 fifo_array_reg_8__19_ ( .D(n1654), .CLK(clk), .Q(fifo_array[291])
         );
  DFFPOSX1 fifo_array_reg_8__18_ ( .D(n1653), .CLK(clk), .Q(fifo_array[290])
         );
  DFFPOSX1 fifo_array_reg_8__17_ ( .D(n1652), .CLK(clk), .Q(fifo_array[289])
         );
  DFFPOSX1 fifo_array_reg_8__16_ ( .D(n1651), .CLK(clk), .Q(fifo_array[288])
         );
  DFFPOSX1 fifo_array_reg_8__15_ ( .D(n1650), .CLK(clk), .Q(fifo_array[287])
         );
  DFFPOSX1 fifo_array_reg_8__14_ ( .D(n1649), .CLK(clk), .Q(fifo_array[286])
         );
  DFFPOSX1 fifo_array_reg_8__13_ ( .D(n1648), .CLK(clk), .Q(fifo_array[285])
         );
  DFFPOSX1 fifo_array_reg_8__12_ ( .D(n1647), .CLK(clk), .Q(fifo_array[284])
         );
  DFFPOSX1 fifo_array_reg_8__11_ ( .D(n1646), .CLK(clk), .Q(fifo_array[283])
         );
  DFFPOSX1 fifo_array_reg_8__10_ ( .D(n1645), .CLK(clk), .Q(fifo_array[282])
         );
  DFFPOSX1 fifo_array_reg_8__9_ ( .D(n1644), .CLK(clk), .Q(fifo_array[281]) );
  DFFPOSX1 fifo_array_reg_8__8_ ( .D(n1643), .CLK(clk), .Q(fifo_array[280]) );
  DFFPOSX1 fifo_array_reg_8__7_ ( .D(n1642), .CLK(clk), .Q(fifo_array[279]) );
  DFFPOSX1 fifo_array_reg_8__6_ ( .D(n1641), .CLK(clk), .Q(fifo_array[278]) );
  DFFPOSX1 fifo_array_reg_8__5_ ( .D(n1640), .CLK(clk), .Q(fifo_array[277]) );
  DFFPOSX1 fifo_array_reg_8__4_ ( .D(n1639), .CLK(clk), .Q(fifo_array[276]) );
  DFFPOSX1 fifo_array_reg_8__3_ ( .D(n1638), .CLK(clk), .Q(fifo_array[275]) );
  DFFPOSX1 fifo_array_reg_8__2_ ( .D(n1637), .CLK(clk), .Q(fifo_array[274]) );
  DFFPOSX1 fifo_array_reg_8__1_ ( .D(n1636), .CLK(clk), .Q(fifo_array[273]) );
  DFFPOSX1 fifo_array_reg_8__0_ ( .D(n1635), .CLK(clk), .Q(fifo_array[272]) );
  DFFPOSX1 fifo_array_reg_7__33_ ( .D(n1634), .CLK(clk), .Q(fifo_array[271])
         );
  DFFPOSX1 fifo_array_reg_7__32_ ( .D(n1633), .CLK(clk), .Q(fifo_array[270])
         );
  DFFPOSX1 fifo_array_reg_7__31_ ( .D(n1632), .CLK(clk), .Q(fifo_array[269])
         );
  DFFPOSX1 fifo_array_reg_7__30_ ( .D(n1631), .CLK(clk), .Q(fifo_array[268])
         );
  DFFPOSX1 fifo_array_reg_7__29_ ( .D(n1630), .CLK(clk), .Q(fifo_array[267])
         );
  DFFPOSX1 fifo_array_reg_7__28_ ( .D(n1629), .CLK(clk), .Q(fifo_array[266])
         );
  DFFPOSX1 fifo_array_reg_7__27_ ( .D(n1628), .CLK(clk), .Q(fifo_array[265])
         );
  DFFPOSX1 fifo_array_reg_7__26_ ( .D(n1627), .CLK(clk), .Q(fifo_array[264])
         );
  DFFPOSX1 fifo_array_reg_7__25_ ( .D(n1626), .CLK(clk), .Q(fifo_array[263])
         );
  DFFPOSX1 fifo_array_reg_7__24_ ( .D(n1625), .CLK(clk), .Q(fifo_array[262])
         );
  DFFPOSX1 fifo_array_reg_7__23_ ( .D(n1624), .CLK(clk), .Q(fifo_array[261])
         );
  DFFPOSX1 fifo_array_reg_7__22_ ( .D(n1623), .CLK(clk), .Q(fifo_array[260])
         );
  DFFPOSX1 fifo_array_reg_7__21_ ( .D(n1622), .CLK(clk), .Q(fifo_array[259])
         );
  DFFPOSX1 fifo_array_reg_7__20_ ( .D(n1621), .CLK(clk), .Q(fifo_array[258])
         );
  DFFPOSX1 fifo_array_reg_7__19_ ( .D(n1620), .CLK(clk), .Q(fifo_array[257])
         );
  DFFPOSX1 fifo_array_reg_7__18_ ( .D(n1619), .CLK(clk), .Q(fifo_array[256])
         );
  DFFPOSX1 fifo_array_reg_7__17_ ( .D(n1618), .CLK(clk), .Q(fifo_array[255])
         );
  DFFPOSX1 fifo_array_reg_7__16_ ( .D(n1617), .CLK(clk), .Q(fifo_array[254])
         );
  DFFPOSX1 fifo_array_reg_7__15_ ( .D(n1616), .CLK(clk), .Q(fifo_array[253])
         );
  DFFPOSX1 fifo_array_reg_7__14_ ( .D(n1615), .CLK(clk), .Q(fifo_array[252])
         );
  DFFPOSX1 fifo_array_reg_7__13_ ( .D(n1614), .CLK(clk), .Q(fifo_array[251])
         );
  DFFPOSX1 fifo_array_reg_7__12_ ( .D(n1613), .CLK(clk), .Q(fifo_array[250])
         );
  DFFPOSX1 fifo_array_reg_7__11_ ( .D(n1612), .CLK(clk), .Q(fifo_array[249])
         );
  DFFPOSX1 fifo_array_reg_7__10_ ( .D(n1611), .CLK(clk), .Q(fifo_array[248])
         );
  DFFPOSX1 fifo_array_reg_7__9_ ( .D(n1610), .CLK(clk), .Q(fifo_array[247]) );
  DFFPOSX1 fifo_array_reg_7__8_ ( .D(n1609), .CLK(clk), .Q(fifo_array[246]) );
  DFFPOSX1 fifo_array_reg_7__7_ ( .D(n1608), .CLK(clk), .Q(fifo_array[245]) );
  DFFPOSX1 fifo_array_reg_7__6_ ( .D(n1607), .CLK(clk), .Q(fifo_array[244]) );
  DFFPOSX1 fifo_array_reg_7__5_ ( .D(n1606), .CLK(clk), .Q(fifo_array[243]) );
  DFFPOSX1 fifo_array_reg_7__4_ ( .D(n1605), .CLK(clk), .Q(fifo_array[242]) );
  DFFPOSX1 fifo_array_reg_7__3_ ( .D(n1604), .CLK(clk), .Q(fifo_array[241]) );
  DFFPOSX1 fifo_array_reg_7__2_ ( .D(n1603), .CLK(clk), .Q(fifo_array[240]) );
  DFFPOSX1 fifo_array_reg_7__1_ ( .D(n1602), .CLK(clk), .Q(fifo_array[239]) );
  DFFPOSX1 fifo_array_reg_7__0_ ( .D(n1601), .CLK(clk), .Q(fifo_array[238]) );
  DFFPOSX1 fifo_array_reg_6__33_ ( .D(n1600), .CLK(clk), .Q(fifo_array[237])
         );
  DFFPOSX1 fifo_array_reg_6__32_ ( .D(n1599), .CLK(clk), .Q(fifo_array[236])
         );
  DFFPOSX1 fifo_array_reg_6__31_ ( .D(n1598), .CLK(clk), .Q(fifo_array[235])
         );
  DFFPOSX1 fifo_array_reg_6__30_ ( .D(n1597), .CLK(clk), .Q(fifo_array[234])
         );
  DFFPOSX1 fifo_array_reg_6__29_ ( .D(n1596), .CLK(clk), .Q(fifo_array[233])
         );
  DFFPOSX1 fifo_array_reg_6__28_ ( .D(n1595), .CLK(clk), .Q(fifo_array[232])
         );
  DFFPOSX1 fifo_array_reg_6__27_ ( .D(n1594), .CLK(clk), .Q(fifo_array[231])
         );
  DFFPOSX1 fifo_array_reg_6__26_ ( .D(n1593), .CLK(clk), .Q(fifo_array[230])
         );
  DFFPOSX1 fifo_array_reg_6__25_ ( .D(n1592), .CLK(clk), .Q(fifo_array[229])
         );
  DFFPOSX1 fifo_array_reg_6__24_ ( .D(n1591), .CLK(clk), .Q(fifo_array[228])
         );
  DFFPOSX1 fifo_array_reg_6__23_ ( .D(n1590), .CLK(clk), .Q(fifo_array[227])
         );
  DFFPOSX1 fifo_array_reg_6__22_ ( .D(n1589), .CLK(clk), .Q(fifo_array[226])
         );
  DFFPOSX1 fifo_array_reg_6__21_ ( .D(n1588), .CLK(clk), .Q(fifo_array[225])
         );
  DFFPOSX1 fifo_array_reg_6__20_ ( .D(n1587), .CLK(clk), .Q(fifo_array[224])
         );
  DFFPOSX1 fifo_array_reg_6__19_ ( .D(n1586), .CLK(clk), .Q(fifo_array[223])
         );
  DFFPOSX1 fifo_array_reg_6__18_ ( .D(n1585), .CLK(clk), .Q(fifo_array[222])
         );
  DFFPOSX1 fifo_array_reg_6__17_ ( .D(n1584), .CLK(clk), .Q(fifo_array[221])
         );
  DFFPOSX1 fifo_array_reg_6__16_ ( .D(n1583), .CLK(clk), .Q(fifo_array[220])
         );
  DFFPOSX1 fifo_array_reg_6__15_ ( .D(n1582), .CLK(clk), .Q(fifo_array[219])
         );
  DFFPOSX1 fifo_array_reg_6__14_ ( .D(n1581), .CLK(clk), .Q(fifo_array[218])
         );
  DFFPOSX1 fifo_array_reg_6__13_ ( .D(n1580), .CLK(clk), .Q(fifo_array[217])
         );
  DFFPOSX1 fifo_array_reg_6__12_ ( .D(n1579), .CLK(clk), .Q(fifo_array[216])
         );
  DFFPOSX1 fifo_array_reg_6__11_ ( .D(n1578), .CLK(clk), .Q(fifo_array[215])
         );
  DFFPOSX1 fifo_array_reg_6__10_ ( .D(n1577), .CLK(clk), .Q(fifo_array[214])
         );
  DFFPOSX1 fifo_array_reg_6__9_ ( .D(n1576), .CLK(clk), .Q(fifo_array[213]) );
  DFFPOSX1 fifo_array_reg_6__8_ ( .D(n1575), .CLK(clk), .Q(fifo_array[212]) );
  DFFPOSX1 fifo_array_reg_6__7_ ( .D(n1574), .CLK(clk), .Q(fifo_array[211]) );
  DFFPOSX1 fifo_array_reg_6__6_ ( .D(n1573), .CLK(clk), .Q(fifo_array[210]) );
  DFFPOSX1 fifo_array_reg_6__5_ ( .D(n1572), .CLK(clk), .Q(fifo_array[209]) );
  DFFPOSX1 fifo_array_reg_6__4_ ( .D(n1571), .CLK(clk), .Q(fifo_array[208]) );
  DFFPOSX1 fifo_array_reg_6__3_ ( .D(n1570), .CLK(clk), .Q(fifo_array[207]) );
  DFFPOSX1 fifo_array_reg_6__2_ ( .D(n1569), .CLK(clk), .Q(fifo_array[206]) );
  DFFPOSX1 fifo_array_reg_6__1_ ( .D(n1568), .CLK(clk), .Q(fifo_array[205]) );
  DFFPOSX1 fifo_array_reg_6__0_ ( .D(n1567), .CLK(clk), .Q(fifo_array[204]) );
  DFFPOSX1 fifo_array_reg_5__33_ ( .D(n1566), .CLK(clk), .Q(fifo_array[203])
         );
  DFFPOSX1 fifo_array_reg_5__32_ ( .D(n1565), .CLK(clk), .Q(fifo_array[202])
         );
  DFFPOSX1 fifo_array_reg_5__31_ ( .D(n1564), .CLK(clk), .Q(fifo_array[201])
         );
  DFFPOSX1 fifo_array_reg_5__30_ ( .D(n1563), .CLK(clk), .Q(fifo_array[200])
         );
  DFFPOSX1 fifo_array_reg_5__29_ ( .D(n1562), .CLK(clk), .Q(fifo_array[199])
         );
  DFFPOSX1 fifo_array_reg_5__28_ ( .D(n1561), .CLK(clk), .Q(fifo_array[198])
         );
  DFFPOSX1 fifo_array_reg_5__27_ ( .D(n1560), .CLK(clk), .Q(fifo_array[197])
         );
  DFFPOSX1 fifo_array_reg_5__26_ ( .D(n1559), .CLK(clk), .Q(fifo_array[196])
         );
  DFFPOSX1 fifo_array_reg_5__25_ ( .D(n1558), .CLK(clk), .Q(fifo_array[195])
         );
  DFFPOSX1 fifo_array_reg_5__24_ ( .D(n1557), .CLK(clk), .Q(fifo_array[194])
         );
  DFFPOSX1 fifo_array_reg_5__23_ ( .D(n1556), .CLK(clk), .Q(fifo_array[193])
         );
  DFFPOSX1 fifo_array_reg_5__22_ ( .D(n1555), .CLK(clk), .Q(fifo_array[192])
         );
  DFFPOSX1 fifo_array_reg_5__21_ ( .D(n1554), .CLK(clk), .Q(fifo_array[191])
         );
  DFFPOSX1 fifo_array_reg_5__20_ ( .D(n1553), .CLK(clk), .Q(fifo_array[190])
         );
  DFFPOSX1 fifo_array_reg_5__19_ ( .D(n1552), .CLK(clk), .Q(fifo_array[189])
         );
  DFFPOSX1 fifo_array_reg_5__18_ ( .D(n1551), .CLK(clk), .Q(fifo_array[188])
         );
  DFFPOSX1 fifo_array_reg_5__17_ ( .D(n1550), .CLK(clk), .Q(fifo_array[187])
         );
  DFFPOSX1 fifo_array_reg_5__16_ ( .D(n1549), .CLK(clk), .Q(fifo_array[186])
         );
  DFFPOSX1 fifo_array_reg_5__15_ ( .D(n1548), .CLK(clk), .Q(fifo_array[185])
         );
  DFFPOSX1 fifo_array_reg_5__14_ ( .D(n1547), .CLK(clk), .Q(fifo_array[184])
         );
  DFFPOSX1 fifo_array_reg_5__13_ ( .D(n1546), .CLK(clk), .Q(fifo_array[183])
         );
  DFFPOSX1 fifo_array_reg_5__12_ ( .D(n1545), .CLK(clk), .Q(fifo_array[182])
         );
  DFFPOSX1 fifo_array_reg_5__11_ ( .D(n1544), .CLK(clk), .Q(fifo_array[181])
         );
  DFFPOSX1 fifo_array_reg_5__10_ ( .D(n1543), .CLK(clk), .Q(fifo_array[180])
         );
  DFFPOSX1 fifo_array_reg_5__9_ ( .D(n1542), .CLK(clk), .Q(fifo_array[179]) );
  DFFPOSX1 fifo_array_reg_5__8_ ( .D(n1541), .CLK(clk), .Q(fifo_array[178]) );
  DFFPOSX1 fifo_array_reg_5__7_ ( .D(n1540), .CLK(clk), .Q(fifo_array[177]) );
  DFFPOSX1 fifo_array_reg_5__6_ ( .D(n1539), .CLK(clk), .Q(fifo_array[176]) );
  DFFPOSX1 fifo_array_reg_5__5_ ( .D(n1538), .CLK(clk), .Q(fifo_array[175]) );
  DFFPOSX1 fifo_array_reg_5__4_ ( .D(n1537), .CLK(clk), .Q(fifo_array[174]) );
  DFFPOSX1 fifo_array_reg_5__3_ ( .D(n1536), .CLK(clk), .Q(fifo_array[173]) );
  DFFPOSX1 fifo_array_reg_5__2_ ( .D(n1535), .CLK(clk), .Q(fifo_array[172]) );
  DFFPOSX1 fifo_array_reg_5__1_ ( .D(n1534), .CLK(clk), .Q(fifo_array[171]) );
  DFFPOSX1 fifo_array_reg_5__0_ ( .D(n1533), .CLK(clk), .Q(fifo_array[170]) );
  DFFPOSX1 fifo_array_reg_4__33_ ( .D(n1532), .CLK(clk), .Q(fifo_array[169])
         );
  DFFPOSX1 fifo_array_reg_4__32_ ( .D(n1531), .CLK(clk), .Q(fifo_array[168])
         );
  DFFPOSX1 fifo_array_reg_4__31_ ( .D(n1530), .CLK(clk), .Q(fifo_array[167])
         );
  DFFPOSX1 fifo_array_reg_4__30_ ( .D(n1529), .CLK(clk), .Q(fifo_array[166])
         );
  DFFPOSX1 fifo_array_reg_4__29_ ( .D(n1528), .CLK(clk), .Q(fifo_array[165])
         );
  DFFPOSX1 fifo_array_reg_4__28_ ( .D(n1527), .CLK(clk), .Q(fifo_array[164])
         );
  DFFPOSX1 fifo_array_reg_4__27_ ( .D(n1526), .CLK(clk), .Q(fifo_array[163])
         );
  DFFPOSX1 fifo_array_reg_4__26_ ( .D(n1525), .CLK(clk), .Q(fifo_array[162])
         );
  DFFPOSX1 fifo_array_reg_4__25_ ( .D(n1524), .CLK(clk), .Q(fifo_array[161])
         );
  DFFPOSX1 fifo_array_reg_4__24_ ( .D(n1523), .CLK(clk), .Q(fifo_array[160])
         );
  DFFPOSX1 fifo_array_reg_4__23_ ( .D(n1522), .CLK(clk), .Q(fifo_array[159])
         );
  DFFPOSX1 fifo_array_reg_4__22_ ( .D(n1521), .CLK(clk), .Q(fifo_array[158])
         );
  DFFPOSX1 fifo_array_reg_4__21_ ( .D(n1520), .CLK(clk), .Q(fifo_array[157])
         );
  DFFPOSX1 fifo_array_reg_4__20_ ( .D(n1519), .CLK(clk), .Q(fifo_array[156])
         );
  DFFPOSX1 fifo_array_reg_4__19_ ( .D(n1518), .CLK(clk), .Q(fifo_array[155])
         );
  DFFPOSX1 fifo_array_reg_4__18_ ( .D(n1517), .CLK(clk), .Q(fifo_array[154])
         );
  DFFPOSX1 fifo_array_reg_4__17_ ( .D(n1516), .CLK(clk), .Q(fifo_array[153])
         );
  DFFPOSX1 fifo_array_reg_4__16_ ( .D(n1515), .CLK(clk), .Q(fifo_array[152])
         );
  DFFPOSX1 fifo_array_reg_4__15_ ( .D(n1514), .CLK(clk), .Q(fifo_array[151])
         );
  DFFPOSX1 fifo_array_reg_4__14_ ( .D(n1513), .CLK(clk), .Q(fifo_array[150])
         );
  DFFPOSX1 fifo_array_reg_4__13_ ( .D(n1512), .CLK(clk), .Q(fifo_array[149])
         );
  DFFPOSX1 fifo_array_reg_4__12_ ( .D(n1511), .CLK(clk), .Q(fifo_array[148])
         );
  DFFPOSX1 fifo_array_reg_4__11_ ( .D(n1510), .CLK(clk), .Q(fifo_array[147])
         );
  DFFPOSX1 fifo_array_reg_4__10_ ( .D(n1509), .CLK(clk), .Q(fifo_array[146])
         );
  DFFPOSX1 fifo_array_reg_4__9_ ( .D(n1508), .CLK(clk), .Q(fifo_array[145]) );
  DFFPOSX1 fifo_array_reg_4__8_ ( .D(n1507), .CLK(clk), .Q(fifo_array[144]) );
  DFFPOSX1 fifo_array_reg_4__7_ ( .D(n1506), .CLK(clk), .Q(fifo_array[143]) );
  DFFPOSX1 fifo_array_reg_4__6_ ( .D(n1505), .CLK(clk), .Q(fifo_array[142]) );
  DFFPOSX1 fifo_array_reg_4__5_ ( .D(n1504), .CLK(clk), .Q(fifo_array[141]) );
  DFFPOSX1 fifo_array_reg_4__4_ ( .D(n1503), .CLK(clk), .Q(fifo_array[140]) );
  DFFPOSX1 fifo_array_reg_4__3_ ( .D(n1502), .CLK(clk), .Q(fifo_array[139]) );
  DFFPOSX1 fifo_array_reg_4__2_ ( .D(n1501), .CLK(clk), .Q(fifo_array[138]) );
  DFFPOSX1 fifo_array_reg_4__1_ ( .D(n1500), .CLK(clk), .Q(fifo_array[137]) );
  DFFPOSX1 fifo_array_reg_4__0_ ( .D(n1499), .CLK(clk), .Q(fifo_array[136]) );
  DFFPOSX1 fifo_array_reg_3__33_ ( .D(n1498), .CLK(clk), .Q(fifo_array[135])
         );
  DFFPOSX1 fifo_array_reg_3__32_ ( .D(n1497), .CLK(clk), .Q(fifo_array[134])
         );
  DFFPOSX1 fifo_array_reg_3__31_ ( .D(n1496), .CLK(clk), .Q(fifo_array[133])
         );
  DFFPOSX1 fifo_array_reg_3__30_ ( .D(n1495), .CLK(clk), .Q(fifo_array[132])
         );
  DFFPOSX1 fifo_array_reg_3__29_ ( .D(n1494), .CLK(clk), .Q(fifo_array[131])
         );
  DFFPOSX1 fifo_array_reg_3__28_ ( .D(n1493), .CLK(clk), .Q(fifo_array[130])
         );
  DFFPOSX1 fifo_array_reg_3__27_ ( .D(n1492), .CLK(clk), .Q(fifo_array[129])
         );
  DFFPOSX1 fifo_array_reg_3__26_ ( .D(n1491), .CLK(clk), .Q(fifo_array[128])
         );
  DFFPOSX1 fifo_array_reg_3__25_ ( .D(n1490), .CLK(clk), .Q(fifo_array[127])
         );
  DFFPOSX1 fifo_array_reg_3__24_ ( .D(n1489), .CLK(clk), .Q(fifo_array[126])
         );
  DFFPOSX1 fifo_array_reg_3__23_ ( .D(n1488), .CLK(clk), .Q(fifo_array[125])
         );
  DFFPOSX1 fifo_array_reg_3__22_ ( .D(n1487), .CLK(clk), .Q(fifo_array[124])
         );
  DFFPOSX1 fifo_array_reg_3__21_ ( .D(n1486), .CLK(clk), .Q(fifo_array[123])
         );
  DFFPOSX1 fifo_array_reg_3__20_ ( .D(n1485), .CLK(clk), .Q(fifo_array[122])
         );
  DFFPOSX1 fifo_array_reg_3__19_ ( .D(n1484), .CLK(clk), .Q(fifo_array[121])
         );
  DFFPOSX1 fifo_array_reg_3__18_ ( .D(n1483), .CLK(clk), .Q(fifo_array[120])
         );
  DFFPOSX1 fifo_array_reg_3__17_ ( .D(n1482), .CLK(clk), .Q(fifo_array[119])
         );
  DFFPOSX1 fifo_array_reg_3__16_ ( .D(n1481), .CLK(clk), .Q(fifo_array[118])
         );
  DFFPOSX1 fifo_array_reg_3__15_ ( .D(n1480), .CLK(clk), .Q(fifo_array[117])
         );
  DFFPOSX1 fifo_array_reg_3__14_ ( .D(n1479), .CLK(clk), .Q(fifo_array[116])
         );
  DFFPOSX1 fifo_array_reg_3__13_ ( .D(n1478), .CLK(clk), .Q(fifo_array[115])
         );
  DFFPOSX1 fifo_array_reg_3__12_ ( .D(n1477), .CLK(clk), .Q(fifo_array[114])
         );
  DFFPOSX1 fifo_array_reg_3__11_ ( .D(n1476), .CLK(clk), .Q(fifo_array[113])
         );
  DFFPOSX1 fifo_array_reg_3__10_ ( .D(n1475), .CLK(clk), .Q(fifo_array[112])
         );
  DFFPOSX1 fifo_array_reg_3__9_ ( .D(n1474), .CLK(clk), .Q(fifo_array[111]) );
  DFFPOSX1 fifo_array_reg_3__8_ ( .D(n1473), .CLK(clk), .Q(fifo_array[110]) );
  DFFPOSX1 fifo_array_reg_3__7_ ( .D(n1472), .CLK(clk), .Q(fifo_array[109]) );
  DFFPOSX1 fifo_array_reg_3__6_ ( .D(n1471), .CLK(clk), .Q(fifo_array[108]) );
  DFFPOSX1 fifo_array_reg_3__5_ ( .D(n1470), .CLK(clk), .Q(fifo_array[107]) );
  DFFPOSX1 fifo_array_reg_3__4_ ( .D(n1469), .CLK(clk), .Q(fifo_array[106]) );
  DFFPOSX1 fifo_array_reg_3__3_ ( .D(n1468), .CLK(clk), .Q(fifo_array[105]) );
  DFFPOSX1 fifo_array_reg_3__2_ ( .D(n1467), .CLK(clk), .Q(fifo_array[104]) );
  DFFPOSX1 fifo_array_reg_3__1_ ( .D(n1466), .CLK(clk), .Q(fifo_array[103]) );
  DFFPOSX1 fifo_array_reg_3__0_ ( .D(n1465), .CLK(clk), .Q(fifo_array[102]) );
  DFFPOSX1 fifo_array_reg_2__33_ ( .D(n1464), .CLK(clk), .Q(fifo_array[101])
         );
  DFFPOSX1 fifo_array_reg_2__32_ ( .D(n1463), .CLK(clk), .Q(fifo_array[100])
         );
  DFFPOSX1 fifo_array_reg_2__31_ ( .D(n1462), .CLK(clk), .Q(fifo_array[99]) );
  DFFPOSX1 fifo_array_reg_2__30_ ( .D(n1461), .CLK(clk), .Q(fifo_array[98]) );
  DFFPOSX1 fifo_array_reg_2__29_ ( .D(n1460), .CLK(clk), .Q(fifo_array[97]) );
  DFFPOSX1 fifo_array_reg_2__28_ ( .D(n1459), .CLK(clk), .Q(fifo_array[96]) );
  DFFPOSX1 fifo_array_reg_2__27_ ( .D(n1458), .CLK(clk), .Q(fifo_array[95]) );
  DFFPOSX1 fifo_array_reg_2__26_ ( .D(n1457), .CLK(clk), .Q(fifo_array[94]) );
  DFFPOSX1 fifo_array_reg_2__25_ ( .D(n1456), .CLK(clk), .Q(fifo_array[93]) );
  DFFPOSX1 fifo_array_reg_2__24_ ( .D(n1455), .CLK(clk), .Q(fifo_array[92]) );
  DFFPOSX1 fifo_array_reg_2__23_ ( .D(n1454), .CLK(clk), .Q(fifo_array[91]) );
  DFFPOSX1 fifo_array_reg_2__22_ ( .D(n1453), .CLK(clk), .Q(fifo_array[90]) );
  DFFPOSX1 fifo_array_reg_2__21_ ( .D(n1452), .CLK(clk), .Q(fifo_array[89]) );
  DFFPOSX1 fifo_array_reg_2__20_ ( .D(n1451), .CLK(clk), .Q(fifo_array[88]) );
  DFFPOSX1 fifo_array_reg_2__19_ ( .D(n1450), .CLK(clk), .Q(fifo_array[87]) );
  DFFPOSX1 fifo_array_reg_2__18_ ( .D(n1449), .CLK(clk), .Q(fifo_array[86]) );
  DFFPOSX1 fifo_array_reg_2__17_ ( .D(n1448), .CLK(clk), .Q(fifo_array[85]) );
  DFFPOSX1 fifo_array_reg_2__16_ ( .D(n1447), .CLK(clk), .Q(fifo_array[84]) );
  DFFPOSX1 fifo_array_reg_2__15_ ( .D(n1446), .CLK(clk), .Q(fifo_array[83]) );
  DFFPOSX1 fifo_array_reg_2__14_ ( .D(n1445), .CLK(clk), .Q(fifo_array[82]) );
  DFFPOSX1 fifo_array_reg_2__13_ ( .D(n1444), .CLK(clk), .Q(fifo_array[81]) );
  DFFPOSX1 fifo_array_reg_2__12_ ( .D(n1443), .CLK(clk), .Q(fifo_array[80]) );
  DFFPOSX1 fifo_array_reg_2__11_ ( .D(n1442), .CLK(clk), .Q(fifo_array[79]) );
  DFFPOSX1 fifo_array_reg_2__10_ ( .D(n1441), .CLK(clk), .Q(fifo_array[78]) );
  DFFPOSX1 fifo_array_reg_2__9_ ( .D(n1440), .CLK(clk), .Q(fifo_array[77]) );
  DFFPOSX1 fifo_array_reg_2__8_ ( .D(n1439), .CLK(clk), .Q(fifo_array[76]) );
  DFFPOSX1 fifo_array_reg_2__7_ ( .D(n1438), .CLK(clk), .Q(fifo_array[75]) );
  DFFPOSX1 fifo_array_reg_2__6_ ( .D(n1437), .CLK(clk), .Q(fifo_array[74]) );
  DFFPOSX1 fifo_array_reg_2__5_ ( .D(n1436), .CLK(clk), .Q(fifo_array[73]) );
  DFFPOSX1 fifo_array_reg_2__4_ ( .D(n1435), .CLK(clk), .Q(fifo_array[72]) );
  DFFPOSX1 fifo_array_reg_2__3_ ( .D(n1434), .CLK(clk), .Q(fifo_array[71]) );
  DFFPOSX1 fifo_array_reg_2__2_ ( .D(n1433), .CLK(clk), .Q(fifo_array[70]) );
  DFFPOSX1 fifo_array_reg_2__1_ ( .D(n1432), .CLK(clk), .Q(fifo_array[69]) );
  DFFPOSX1 fifo_array_reg_2__0_ ( .D(n1431), .CLK(clk), .Q(fifo_array[68]) );
  DFFPOSX1 fifo_array_reg_1__33_ ( .D(n1430), .CLK(clk), .Q(fifo_array[67]) );
  DFFPOSX1 fifo_array_reg_1__32_ ( .D(n1429), .CLK(clk), .Q(fifo_array[66]) );
  DFFPOSX1 fifo_array_reg_1__31_ ( .D(n1428), .CLK(clk), .Q(fifo_array[65]) );
  DFFPOSX1 fifo_array_reg_1__30_ ( .D(n1427), .CLK(clk), .Q(fifo_array[64]) );
  DFFPOSX1 fifo_array_reg_1__29_ ( .D(n1426), .CLK(clk), .Q(fifo_array[63]) );
  DFFPOSX1 fifo_array_reg_1__28_ ( .D(n1425), .CLK(clk), .Q(fifo_array[62]) );
  DFFPOSX1 fifo_array_reg_1__27_ ( .D(n1424), .CLK(clk), .Q(fifo_array[61]) );
  DFFPOSX1 fifo_array_reg_1__26_ ( .D(n1423), .CLK(clk), .Q(fifo_array[60]) );
  DFFPOSX1 fifo_array_reg_1__25_ ( .D(n1422), .CLK(clk), .Q(fifo_array[59]) );
  DFFPOSX1 fifo_array_reg_1__24_ ( .D(n1421), .CLK(clk), .Q(fifo_array[58]) );
  DFFPOSX1 fifo_array_reg_1__23_ ( .D(n1420), .CLK(clk), .Q(fifo_array[57]) );
  DFFPOSX1 fifo_array_reg_1__22_ ( .D(n1419), .CLK(clk), .Q(fifo_array[56]) );
  DFFPOSX1 fifo_array_reg_1__21_ ( .D(n1418), .CLK(clk), .Q(fifo_array[55]) );
  DFFPOSX1 fifo_array_reg_1__20_ ( .D(n1417), .CLK(clk), .Q(fifo_array[54]) );
  DFFPOSX1 fifo_array_reg_1__19_ ( .D(n1416), .CLK(clk), .Q(fifo_array[53]) );
  DFFPOSX1 fifo_array_reg_1__18_ ( .D(n1415), .CLK(clk), .Q(fifo_array[52]) );
  DFFPOSX1 fifo_array_reg_1__17_ ( .D(n1414), .CLK(clk), .Q(fifo_array[51]) );
  DFFPOSX1 fifo_array_reg_1__16_ ( .D(n1413), .CLK(clk), .Q(fifo_array[50]) );
  DFFPOSX1 fifo_array_reg_1__15_ ( .D(n1412), .CLK(clk), .Q(fifo_array[49]) );
  DFFPOSX1 fifo_array_reg_1__14_ ( .D(n1411), .CLK(clk), .Q(fifo_array[48]) );
  DFFPOSX1 fifo_array_reg_1__13_ ( .D(n1410), .CLK(clk), .Q(fifo_array[47]) );
  DFFPOSX1 fifo_array_reg_1__12_ ( .D(n1409), .CLK(clk), .Q(fifo_array[46]) );
  DFFPOSX1 fifo_array_reg_1__11_ ( .D(n1408), .CLK(clk), .Q(fifo_array[45]) );
  DFFPOSX1 fifo_array_reg_1__10_ ( .D(n1407), .CLK(clk), .Q(fifo_array[44]) );
  DFFPOSX1 fifo_array_reg_1__9_ ( .D(n1406), .CLK(clk), .Q(fifo_array[43]) );
  DFFPOSX1 fifo_array_reg_1__8_ ( .D(n1405), .CLK(clk), .Q(fifo_array[42]) );
  DFFPOSX1 fifo_array_reg_1__7_ ( .D(n1404), .CLK(clk), .Q(fifo_array[41]) );
  DFFPOSX1 fifo_array_reg_1__6_ ( .D(n1403), .CLK(clk), .Q(fifo_array[40]) );
  DFFPOSX1 fifo_array_reg_1__5_ ( .D(n1402), .CLK(clk), .Q(fifo_array[39]) );
  DFFPOSX1 fifo_array_reg_1__4_ ( .D(n1401), .CLK(clk), .Q(fifo_array[38]) );
  DFFPOSX1 fifo_array_reg_1__3_ ( .D(n1400), .CLK(clk), .Q(fifo_array[37]) );
  DFFPOSX1 fifo_array_reg_1__2_ ( .D(n1399), .CLK(clk), .Q(fifo_array[36]) );
  DFFPOSX1 fifo_array_reg_1__1_ ( .D(n1398), .CLK(clk), .Q(fifo_array[35]) );
  DFFPOSX1 fifo_array_reg_1__0_ ( .D(n1397), .CLK(clk), .Q(fifo_array[34]) );
  DFFPOSX1 fifo_array_reg_0__33_ ( .D(n1396), .CLK(clk), .Q(fifo_array[33]) );
  DFFPOSX1 fifo_array_reg_0__32_ ( .D(n1395), .CLK(clk), .Q(fifo_array[32]) );
  DFFPOSX1 fifo_array_reg_0__31_ ( .D(n1394), .CLK(clk), .Q(fifo_array[31]) );
  DFFPOSX1 fifo_array_reg_0__30_ ( .D(n1393), .CLK(clk), .Q(fifo_array[30]) );
  DFFPOSX1 fifo_array_reg_0__29_ ( .D(n1392), .CLK(clk), .Q(fifo_array[29]) );
  DFFPOSX1 fifo_array_reg_0__28_ ( .D(n1391), .CLK(clk), .Q(fifo_array[28]) );
  DFFPOSX1 fifo_array_reg_0__27_ ( .D(n1390), .CLK(clk), .Q(fifo_array[27]) );
  DFFPOSX1 fifo_array_reg_0__26_ ( .D(n1389), .CLK(clk), .Q(fifo_array[26]) );
  DFFPOSX1 fifo_array_reg_0__25_ ( .D(n1388), .CLK(clk), .Q(fifo_array[25]) );
  DFFPOSX1 fifo_array_reg_0__24_ ( .D(n1387), .CLK(clk), .Q(fifo_array[24]) );
  DFFPOSX1 fifo_array_reg_0__23_ ( .D(n1386), .CLK(clk), .Q(fifo_array[23]) );
  DFFPOSX1 fifo_array_reg_0__22_ ( .D(n1385), .CLK(clk), .Q(fifo_array[22]) );
  DFFPOSX1 fifo_array_reg_0__21_ ( .D(n1384), .CLK(clk), .Q(fifo_array[21]) );
  DFFPOSX1 fifo_array_reg_0__20_ ( .D(n1383), .CLK(clk), .Q(fifo_array[20]) );
  DFFPOSX1 fifo_array_reg_0__19_ ( .D(n1382), .CLK(clk), .Q(fifo_array[19]) );
  DFFPOSX1 fifo_array_reg_0__18_ ( .D(n1381), .CLK(clk), .Q(fifo_array[18]) );
  DFFPOSX1 fifo_array_reg_0__17_ ( .D(n1380), .CLK(clk), .Q(fifo_array[17]) );
  DFFPOSX1 fifo_array_reg_0__16_ ( .D(n1379), .CLK(clk), .Q(fifo_array[16]) );
  DFFPOSX1 fifo_array_reg_0__15_ ( .D(n1378), .CLK(clk), .Q(fifo_array[15]) );
  DFFPOSX1 fifo_array_reg_0__14_ ( .D(n1377), .CLK(clk), .Q(fifo_array[14]) );
  DFFPOSX1 fifo_array_reg_0__13_ ( .D(n1376), .CLK(clk), .Q(fifo_array[13]) );
  DFFPOSX1 fifo_array_reg_0__12_ ( .D(n1375), .CLK(clk), .Q(fifo_array[12]) );
  DFFPOSX1 fifo_array_reg_0__11_ ( .D(n1374), .CLK(clk), .Q(fifo_array[11]) );
  DFFPOSX1 fifo_array_reg_0__10_ ( .D(n1373), .CLK(clk), .Q(fifo_array[10]) );
  DFFPOSX1 fifo_array_reg_0__9_ ( .D(n1372), .CLK(clk), .Q(fifo_array[9]) );
  DFFPOSX1 fifo_array_reg_0__8_ ( .D(n1371), .CLK(clk), .Q(fifo_array[8]) );
  DFFPOSX1 fifo_array_reg_0__7_ ( .D(n1370), .CLK(clk), .Q(fifo_array[7]) );
  DFFPOSX1 fifo_array_reg_0__6_ ( .D(n1369), .CLK(clk), .Q(fifo_array[6]) );
  DFFPOSX1 fifo_array_reg_0__5_ ( .D(n1368), .CLK(clk), .Q(fifo_array[5]) );
  DFFPOSX1 fifo_array_reg_0__4_ ( .D(n1367), .CLK(clk), .Q(fifo_array[4]) );
  DFFPOSX1 fifo_array_reg_0__3_ ( .D(n1366), .CLK(clk), .Q(fifo_array[3]) );
  DFFPOSX1 fifo_array_reg_0__2_ ( .D(n1365), .CLK(clk), .Q(fifo_array[2]) );
  DFFPOSX1 fifo_array_reg_0__1_ ( .D(n1364), .CLK(clk), .Q(fifo_array[1]) );
  DFFPOSX1 fifo_array_reg_0__0_ ( .D(n1363), .CLK(clk), .Q(fifo_array[0]) );
  OAI21X1 U103 ( .A(n4757), .B(n4664), .C(n3519), .Y(n1363) );
  OAI21X1 U105 ( .A(n4756), .B(n4663), .C(n3452), .Y(n1364) );
  OAI21X1 U107 ( .A(n4756), .B(n4662), .C(n3387), .Y(n1365) );
  OAI21X1 U109 ( .A(n4756), .B(n4661), .C(n3321), .Y(n1366) );
  OAI21X1 U111 ( .A(n4756), .B(n4660), .C(n3253), .Y(n1367) );
  OAI21X1 U113 ( .A(n4756), .B(n4690), .C(n3195), .Y(n1368) );
  OAI21X1 U115 ( .A(n4756), .B(n4689), .C(n3138), .Y(n1369) );
  OAI21X1 U117 ( .A(n4756), .B(n4688), .C(n3080), .Y(n1370) );
  OAI21X1 U119 ( .A(n4756), .B(n4687), .C(n3022), .Y(n1371) );
  OAI21X1 U121 ( .A(n4756), .B(n4686), .C(n3518), .Y(n1372) );
  OAI21X1 U123 ( .A(n4756), .B(n4685), .C(n2968), .Y(n1373) );
  OAI21X1 U125 ( .A(n4756), .B(n4684), .C(n2914), .Y(n1374) );
  OAI21X1 U127 ( .A(n4756), .B(n4683), .C(n2860), .Y(n1375) );
  OAI21X1 U129 ( .A(n4757), .B(n4682), .C(n3451), .Y(n1376) );
  OAI21X1 U131 ( .A(n4756), .B(n4681), .C(n3386), .Y(n1377) );
  OAI21X1 U133 ( .A(n4757), .B(n4680), .C(n3320), .Y(n1378) );
  OAI21X1 U135 ( .A(n4756), .B(n4679), .C(n3252), .Y(n1379) );
  OAI21X1 U137 ( .A(n4757), .B(n4678), .C(n3194), .Y(n1380) );
  OAI21X1 U139 ( .A(n4756), .B(n4677), .C(n3137), .Y(n1381) );
  OAI21X1 U141 ( .A(n4757), .B(n4676), .C(n3079), .Y(n1382) );
  OAI21X1 U143 ( .A(n4756), .B(n4675), .C(n3021), .Y(n1383) );
  OAI21X1 U145 ( .A(n4757), .B(n4674), .C(n2967), .Y(n1384) );
  OAI21X1 U147 ( .A(n4756), .B(n4673), .C(n2913), .Y(n1385) );
  OAI21X1 U149 ( .A(n4757), .B(n4672), .C(n2806), .Y(n1386) );
  OAI21X1 U151 ( .A(n4756), .B(n4671), .C(n2754), .Y(n1387) );
  OAI21X1 U153 ( .A(n4756), .B(n4670), .C(n2702), .Y(n1388) );
  OAI21X1 U155 ( .A(n4756), .B(n4669), .C(n2650), .Y(n1389) );
  OAI21X1 U157 ( .A(n4757), .B(n4668), .C(n2598), .Y(n1390) );
  OAI21X1 U159 ( .A(n4756), .B(n4667), .C(n2597), .Y(n1391) );
  OAI21X1 U161 ( .A(n4756), .B(n4666), .C(n2859), .Y(n1392) );
  OAI21X1 U163 ( .A(n4756), .B(n4665), .C(n2596), .Y(n1393) );
  OAI21X1 U165 ( .A(n4756), .B(n4659), .C(n2595), .Y(n1394) );
  OAI21X1 U167 ( .A(n4756), .B(n4658), .C(n2594), .Y(n1395) );
  OAI21X1 U169 ( .A(n4756), .B(n4657), .C(n2593), .Y(n1396) );
  OAI21X1 U172 ( .A(n4664), .B(n4754), .C(n3450), .Y(n1397) );
  OAI21X1 U174 ( .A(n4663), .B(n4754), .C(n3517), .Y(n1398) );
  OAI21X1 U176 ( .A(n4662), .B(n4754), .C(n3319), .Y(n1399) );
  OAI21X1 U178 ( .A(n4661), .B(n4754), .C(n3385), .Y(n1400) );
  OAI21X1 U180 ( .A(n4660), .B(n4754), .C(n3193), .Y(n1401) );
  OAI21X1 U182 ( .A(n4690), .B(n4754), .C(n3251), .Y(n1402) );
  OAI21X1 U184 ( .A(n4689), .B(n4754), .C(n3078), .Y(n1403) );
  OAI21X1 U186 ( .A(n4688), .B(n4754), .C(n3136), .Y(n1404) );
  OAI21X1 U188 ( .A(n4687), .B(n4754), .C(n2966), .Y(n1405) );
  OAI21X1 U190 ( .A(n4686), .B(n4754), .C(n3449), .Y(n1406) );
  OAI21X1 U192 ( .A(n4685), .B(n4754), .C(n3020), .Y(n1407) );
  OAI21X1 U194 ( .A(n4684), .B(n4754), .C(n2858), .Y(n1408) );
  OAI21X1 U196 ( .A(n4683), .B(n4754), .C(n2912), .Y(n1409) );
  OAI21X1 U198 ( .A(n4682), .B(n4754), .C(n3516), .Y(n1410) );
  OAI21X1 U200 ( .A(n4681), .B(n4755), .C(n3318), .Y(n1411) );
  OAI21X1 U202 ( .A(n4680), .B(n4754), .C(n3384), .Y(n1412) );
  OAI21X1 U204 ( .A(n4679), .B(n4755), .C(n3192), .Y(n1413) );
  OAI21X1 U206 ( .A(n4678), .B(n4754), .C(n3250), .Y(n1414) );
  OAI21X1 U208 ( .A(n4677), .B(n4755), .C(n3077), .Y(n1415) );
  OAI21X1 U210 ( .A(n4676), .B(n4754), .C(n3135), .Y(n1416) );
  OAI21X1 U212 ( .A(n4675), .B(n4755), .C(n2965), .Y(n1417) );
  OAI21X1 U214 ( .A(n4674), .B(n4754), .C(n3019), .Y(n1418) );
  OAI21X1 U216 ( .A(n4673), .B(n4755), .C(n2857), .Y(n1419) );
  OAI21X1 U218 ( .A(n4672), .B(n4754), .C(n2753), .Y(n1420) );
  OAI21X1 U220 ( .A(n4671), .B(n4754), .C(n2805), .Y(n1421) );
  OAI21X1 U222 ( .A(n4670), .B(n4754), .C(n2649), .Y(n1422) );
  OAI21X1 U224 ( .A(n4669), .B(n4754), .C(n2701), .Y(n1423) );
  OAI21X1 U226 ( .A(n4668), .B(n4754), .C(n2592), .Y(n1424) );
  OAI21X1 U228 ( .A(n4667), .B(n4754), .C(n2591), .Y(n1425) );
  OAI21X1 U230 ( .A(n4666), .B(n4755), .C(n2911), .Y(n1426) );
  OAI21X1 U232 ( .A(n4665), .B(n4754), .C(n2590), .Y(n1427) );
  OAI21X1 U234 ( .A(n4659), .B(n4754), .C(n2589), .Y(n1428) );
  OAI21X1 U236 ( .A(n4658), .B(n4754), .C(n2588), .Y(n1429) );
  OAI21X1 U238 ( .A(n4657), .B(n4754), .C(n2587), .Y(n1430) );
  OAI21X1 U241 ( .A(n4664), .B(n4752), .C(n3383), .Y(n1431) );
  OAI21X1 U243 ( .A(n4663), .B(n4752), .C(n3317), .Y(n1432) );
  OAI21X1 U245 ( .A(n4662), .B(n4752), .C(n3515), .Y(n1433) );
  OAI21X1 U247 ( .A(n4661), .B(n4752), .C(n3448), .Y(n1434) );
  OAI21X1 U249 ( .A(n4660), .B(n4752), .C(n3134), .Y(n1435) );
  OAI21X1 U251 ( .A(n4690), .B(n4752), .C(n3076), .Y(n1436) );
  OAI21X1 U253 ( .A(n4689), .B(n4752), .C(n3249), .Y(n1437) );
  OAI21X1 U255 ( .A(n4688), .B(n4752), .C(n3191), .Y(n1438) );
  OAI21X1 U257 ( .A(n4687), .B(n4752), .C(n2910), .Y(n1439) );
  OAI21X1 U259 ( .A(n4686), .B(n4752), .C(n3382), .Y(n1440) );
  OAI21X1 U261 ( .A(n4685), .B(n4752), .C(n2856), .Y(n1441) );
  OAI21X1 U263 ( .A(n4684), .B(n4752), .C(n3018), .Y(n1442) );
  OAI21X1 U265 ( .A(n4683), .B(n4752), .C(n2964), .Y(n1443) );
  OAI21X1 U267 ( .A(n4682), .B(n4752), .C(n3316), .Y(n1444) );
  OAI21X1 U269 ( .A(n4681), .B(n4753), .C(n3514), .Y(n1445) );
  OAI21X1 U271 ( .A(n4680), .B(n4752), .C(n3447), .Y(n1446) );
  OAI21X1 U273 ( .A(n4679), .B(n4753), .C(n3133), .Y(n1447) );
  OAI21X1 U275 ( .A(n4678), .B(n4752), .C(n3075), .Y(n1448) );
  OAI21X1 U277 ( .A(n4677), .B(n4753), .C(n3248), .Y(n1449) );
  OAI21X1 U279 ( .A(n4676), .B(n4752), .C(n3190), .Y(n1450) );
  OAI21X1 U281 ( .A(n4675), .B(n4753), .C(n2909), .Y(n1451) );
  OAI21X1 U283 ( .A(n4674), .B(n4752), .C(n2855), .Y(n1452) );
  OAI21X1 U285 ( .A(n4673), .B(n4753), .C(n3017), .Y(n1453) );
  OAI21X1 U287 ( .A(n4672), .B(n4752), .C(n2700), .Y(n1454) );
  OAI21X1 U289 ( .A(n4671), .B(n4752), .C(n2648), .Y(n1455) );
  OAI21X1 U291 ( .A(n4670), .B(n4752), .C(n2804), .Y(n1456) );
  OAI21X1 U293 ( .A(n4669), .B(n4752), .C(n2752), .Y(n1457) );
  OAI21X1 U295 ( .A(n4668), .B(n4752), .C(n2586), .Y(n1458) );
  OAI21X1 U297 ( .A(n4667), .B(n4752), .C(n2585), .Y(n1459) );
  OAI21X1 U299 ( .A(n4666), .B(n4753), .C(n2963), .Y(n1460) );
  OAI21X1 U301 ( .A(n4665), .B(n4752), .C(n2584), .Y(n1461) );
  OAI21X1 U303 ( .A(n4659), .B(n4752), .C(n2583), .Y(n1462) );
  OAI21X1 U305 ( .A(n4658), .B(n4752), .C(n2582), .Y(n1463) );
  OAI21X1 U307 ( .A(n4657), .B(n4752), .C(n2581), .Y(n1464) );
  OAI21X1 U310 ( .A(n4664), .B(n4750), .C(n3315), .Y(n1465) );
  OAI21X1 U312 ( .A(n4663), .B(n4750), .C(n3381), .Y(n1466) );
  OAI21X1 U314 ( .A(n4662), .B(n4750), .C(n3446), .Y(n1467) );
  OAI21X1 U316 ( .A(n4661), .B(n4750), .C(n3513), .Y(n1468) );
  OAI21X1 U318 ( .A(n4660), .B(n4750), .C(n3074), .Y(n1469) );
  OAI21X1 U320 ( .A(n4690), .B(n4750), .C(n3132), .Y(n1470) );
  OAI21X1 U322 ( .A(n4689), .B(n4750), .C(n3189), .Y(n1471) );
  OAI21X1 U324 ( .A(n4688), .B(n4750), .C(n3247), .Y(n1472) );
  OAI21X1 U326 ( .A(n4687), .B(n4750), .C(n2854), .Y(n1473) );
  OAI21X1 U328 ( .A(n4686), .B(n4750), .C(n3314), .Y(n1474) );
  OAI21X1 U330 ( .A(n4685), .B(n4750), .C(n2908), .Y(n1475) );
  OAI21X1 U332 ( .A(n4684), .B(n4750), .C(n2962), .Y(n1476) );
  OAI21X1 U334 ( .A(n4683), .B(n4750), .C(n3016), .Y(n1477) );
  OAI21X1 U336 ( .A(n4682), .B(n4750), .C(n3380), .Y(n1478) );
  OAI21X1 U338 ( .A(n4681), .B(n4751), .C(n3445), .Y(n1479) );
  OAI21X1 U340 ( .A(n4680), .B(n4750), .C(n3512), .Y(n1480) );
  OAI21X1 U342 ( .A(n4679), .B(n4751), .C(n3073), .Y(n1481) );
  OAI21X1 U344 ( .A(n4678), .B(n4750), .C(n3131), .Y(n1482) );
  OAI21X1 U346 ( .A(n4677), .B(n4751), .C(n3188), .Y(n1483) );
  OAI21X1 U348 ( .A(n4676), .B(n4750), .C(n3246), .Y(n1484) );
  OAI21X1 U350 ( .A(n4675), .B(n4751), .C(n2853), .Y(n1485) );
  OAI21X1 U352 ( .A(n4674), .B(n4750), .C(n2907), .Y(n1486) );
  OAI21X1 U354 ( .A(n4673), .B(n4751), .C(n2961), .Y(n1487) );
  OAI21X1 U356 ( .A(n4672), .B(n4750), .C(n2647), .Y(n1488) );
  OAI21X1 U358 ( .A(n4671), .B(n4750), .C(n2699), .Y(n1489) );
  OAI21X1 U360 ( .A(n4670), .B(n4750), .C(n2751), .Y(n1490) );
  OAI21X1 U362 ( .A(n4669), .B(n4750), .C(n2803), .Y(n1491) );
  OAI21X1 U364 ( .A(n4668), .B(n4750), .C(n2580), .Y(n1492) );
  OAI21X1 U366 ( .A(n4667), .B(n4750), .C(n2579), .Y(n1493) );
  OAI21X1 U368 ( .A(n4666), .B(n4751), .C(n3015), .Y(n1494) );
  OAI21X1 U370 ( .A(n4665), .B(n4750), .C(n2578), .Y(n1495) );
  OAI21X1 U372 ( .A(n4659), .B(n4750), .C(n2577), .Y(n1496) );
  OAI21X1 U374 ( .A(n4658), .B(n4750), .C(n2576), .Y(n1497) );
  OAI21X1 U376 ( .A(n4657), .B(n4750), .C(n2575), .Y(n1498) );
  OAI21X1 U379 ( .A(n4664), .B(n4748), .C(n3245), .Y(n1499) );
  OAI21X1 U381 ( .A(n4663), .B(n4748), .C(n3187), .Y(n1500) );
  OAI21X1 U383 ( .A(n4662), .B(n4748), .C(n3130), .Y(n1501) );
  OAI21X1 U385 ( .A(n4661), .B(n4748), .C(n3072), .Y(n1502) );
  OAI21X1 U387 ( .A(n4660), .B(n4748), .C(n3511), .Y(n1503) );
  OAI21X1 U389 ( .A(n4690), .B(n4748), .C(n3444), .Y(n1504) );
  OAI21X1 U391 ( .A(n4689), .B(n4748), .C(n3379), .Y(n1505) );
  OAI21X1 U393 ( .A(n4688), .B(n4748), .C(n3313), .Y(n1506) );
  OAI21X1 U395 ( .A(n4687), .B(n4748), .C(n2802), .Y(n1507) );
  OAI21X1 U397 ( .A(n4686), .B(n4748), .C(n3244), .Y(n1508) );
  OAI21X1 U399 ( .A(n4685), .B(n4748), .C(n2750), .Y(n1509) );
  OAI21X1 U401 ( .A(n4684), .B(n4748), .C(n2698), .Y(n1510) );
  OAI21X1 U403 ( .A(n4683), .B(n4748), .C(n2646), .Y(n1511) );
  OAI21X1 U405 ( .A(n4682), .B(n4748), .C(n3186), .Y(n1512) );
  OAI21X1 U407 ( .A(n4681), .B(n4749), .C(n3129), .Y(n1513) );
  OAI21X1 U409 ( .A(n4680), .B(n4748), .C(n3071), .Y(n1514) );
  OAI21X1 U411 ( .A(n4679), .B(n4749), .C(n3510), .Y(n1515) );
  OAI21X1 U413 ( .A(n4678), .B(n4748), .C(n3443), .Y(n1516) );
  OAI21X1 U415 ( .A(n4677), .B(n4749), .C(n3378), .Y(n1517) );
  OAI21X1 U417 ( .A(n4676), .B(n4748), .C(n3312), .Y(n1518) );
  OAI21X1 U419 ( .A(n4675), .B(n4749), .C(n2801), .Y(n1519) );
  OAI21X1 U421 ( .A(n4674), .B(n4748), .C(n2749), .Y(n1520) );
  OAI21X1 U423 ( .A(n4673), .B(n4749), .C(n2697), .Y(n1521) );
  OAI21X1 U425 ( .A(n4672), .B(n4748), .C(n3014), .Y(n1522) );
  OAI21X1 U427 ( .A(n4671), .B(n4748), .C(n2960), .Y(n1523) );
  OAI21X1 U429 ( .A(n4670), .B(n4748), .C(n2906), .Y(n1524) );
  OAI21X1 U431 ( .A(n4669), .B(n4748), .C(n2852), .Y(n1525) );
  OAI21X1 U433 ( .A(n4668), .B(n4748), .C(n2574), .Y(n1526) );
  OAI21X1 U435 ( .A(n4667), .B(n4748), .C(n2573), .Y(n1527) );
  OAI21X1 U437 ( .A(n4666), .B(n4749), .C(n2645), .Y(n1528) );
  OAI21X1 U439 ( .A(n4665), .B(n4748), .C(n2572), .Y(n1529) );
  OAI21X1 U441 ( .A(n4659), .B(n4748), .C(n2571), .Y(n1530) );
  OAI21X1 U443 ( .A(n4658), .B(n4748), .C(n2570), .Y(n1531) );
  OAI21X1 U445 ( .A(n4657), .B(n4748), .C(n2569), .Y(n1532) );
  OAI21X1 U448 ( .A(n4664), .B(n4746), .C(n3185), .Y(n1533) );
  OAI21X1 U450 ( .A(n4663), .B(n4746), .C(n3243), .Y(n1534) );
  OAI21X1 U452 ( .A(n4662), .B(n4746), .C(n3070), .Y(n1535) );
  OAI21X1 U454 ( .A(n4661), .B(n4746), .C(n3128), .Y(n1536) );
  OAI21X1 U456 ( .A(n4660), .B(n4746), .C(n3442), .Y(n1537) );
  OAI21X1 U458 ( .A(n4690), .B(n4746), .C(n3509), .Y(n1538) );
  OAI21X1 U460 ( .A(n4689), .B(n4746), .C(n3311), .Y(n1539) );
  OAI21X1 U462 ( .A(n4688), .B(n4746), .C(n3377), .Y(n1540) );
  OAI21X1 U464 ( .A(n4687), .B(n4746), .C(n2748), .Y(n1541) );
  OAI21X1 U466 ( .A(n4686), .B(n4746), .C(n3184), .Y(n1542) );
  OAI21X1 U468 ( .A(n4685), .B(n4746), .C(n2800), .Y(n1543) );
  OAI21X1 U470 ( .A(n4684), .B(n4746), .C(n2644), .Y(n1544) );
  OAI21X1 U472 ( .A(n4683), .B(n4746), .C(n2696), .Y(n1545) );
  OAI21X1 U474 ( .A(n4682), .B(n4746), .C(n3242), .Y(n1546) );
  OAI21X1 U476 ( .A(n4681), .B(n4747), .C(n3069), .Y(n1547) );
  OAI21X1 U478 ( .A(n4680), .B(n4746), .C(n3127), .Y(n1548) );
  OAI21X1 U480 ( .A(n4679), .B(n4747), .C(n3441), .Y(n1549) );
  OAI21X1 U482 ( .A(n4678), .B(n4746), .C(n3508), .Y(n1550) );
  OAI21X1 U484 ( .A(n4677), .B(n4747), .C(n3310), .Y(n1551) );
  OAI21X1 U486 ( .A(n4676), .B(n4746), .C(n3376), .Y(n1552) );
  OAI21X1 U488 ( .A(n4675), .B(n4747), .C(n2747), .Y(n1553) );
  OAI21X1 U490 ( .A(n4674), .B(n4746), .C(n2799), .Y(n1554) );
  OAI21X1 U492 ( .A(n4673), .B(n4747), .C(n2643), .Y(n1555) );
  OAI21X1 U494 ( .A(n4672), .B(n4746), .C(n2959), .Y(n1556) );
  OAI21X1 U496 ( .A(n4671), .B(n4746), .C(n3013), .Y(n1557) );
  OAI21X1 U498 ( .A(n4670), .B(n4746), .C(n2851), .Y(n1558) );
  OAI21X1 U500 ( .A(n4669), .B(n4746), .C(n2905), .Y(n1559) );
  OAI21X1 U502 ( .A(n4668), .B(n4746), .C(n2568), .Y(n1560) );
  OAI21X1 U504 ( .A(n4667), .B(n4746), .C(n2567), .Y(n1561) );
  OAI21X1 U506 ( .A(n4666), .B(n4747), .C(n2695), .Y(n1562) );
  OAI21X1 U508 ( .A(n4665), .B(n4746), .C(n2566), .Y(n1563) );
  OAI21X1 U510 ( .A(n4659), .B(n4746), .C(n2565), .Y(n1564) );
  OAI21X1 U512 ( .A(n4658), .B(n4746), .C(n2564), .Y(n1565) );
  OAI21X1 U514 ( .A(n4657), .B(n4746), .C(n2563), .Y(n1566) );
  OAI21X1 U517 ( .A(n4664), .B(n4744), .C(n3126), .Y(n1567) );
  OAI21X1 U519 ( .A(n4663), .B(n4744), .C(n3068), .Y(n1568) );
  OAI21X1 U521 ( .A(n4662), .B(n4744), .C(n3241), .Y(n1569) );
  OAI21X1 U523 ( .A(n4661), .B(n4744), .C(n3183), .Y(n1570) );
  OAI21X1 U525 ( .A(n4660), .B(n4744), .C(n3375), .Y(n1571) );
  OAI21X1 U527 ( .A(n4690), .B(n4744), .C(n3309), .Y(n1572) );
  OAI21X1 U529 ( .A(n4689), .B(n4744), .C(n3507), .Y(n1573) );
  OAI21X1 U531 ( .A(n4688), .B(n4744), .C(n3440), .Y(n1574) );
  OAI21X1 U533 ( .A(n4687), .B(n4744), .C(n2694), .Y(n1575) );
  OAI21X1 U535 ( .A(n4686), .B(n4744), .C(n3125), .Y(n1576) );
  OAI21X1 U537 ( .A(n4685), .B(n4744), .C(n2642), .Y(n1577) );
  OAI21X1 U539 ( .A(n4684), .B(n4744), .C(n2798), .Y(n1578) );
  OAI21X1 U541 ( .A(n4683), .B(n4744), .C(n2746), .Y(n1579) );
  OAI21X1 U543 ( .A(n4682), .B(n4744), .C(n3067), .Y(n1580) );
  OAI21X1 U545 ( .A(n4681), .B(n4745), .C(n3240), .Y(n1581) );
  OAI21X1 U547 ( .A(n4680), .B(n4744), .C(n3182), .Y(n1582) );
  OAI21X1 U549 ( .A(n4679), .B(n4745), .C(n3374), .Y(n1583) );
  OAI21X1 U551 ( .A(n4678), .B(n4744), .C(n3308), .Y(n1584) );
  OAI21X1 U553 ( .A(n4677), .B(n4745), .C(n3506), .Y(n1585) );
  OAI21X1 U555 ( .A(n4676), .B(n4744), .C(n3439), .Y(n1586) );
  OAI21X1 U557 ( .A(n4675), .B(n4745), .C(n2693), .Y(n1587) );
  OAI21X1 U559 ( .A(n4674), .B(n4744), .C(n2641), .Y(n1588) );
  OAI21X1 U561 ( .A(n4673), .B(n4745), .C(n2797), .Y(n1589) );
  OAI21X1 U563 ( .A(n4672), .B(n4744), .C(n2904), .Y(n1590) );
  OAI21X1 U565 ( .A(n4671), .B(n4744), .C(n2850), .Y(n1591) );
  OAI21X1 U567 ( .A(n4670), .B(n4744), .C(n3012), .Y(n1592) );
  OAI21X1 U569 ( .A(n4669), .B(n4744), .C(n2958), .Y(n1593) );
  OAI21X1 U571 ( .A(n4668), .B(n4744), .C(n2562), .Y(n1594) );
  OAI21X1 U573 ( .A(n4667), .B(n4744), .C(n2561), .Y(n1595) );
  OAI21X1 U575 ( .A(n4666), .B(n4745), .C(n2745), .Y(n1596) );
  OAI21X1 U577 ( .A(n4665), .B(n4744), .C(n2560), .Y(n1597) );
  OAI21X1 U579 ( .A(n4659), .B(n4744), .C(n2559), .Y(n1598) );
  OAI21X1 U581 ( .A(n4658), .B(n4744), .C(n2558), .Y(n1599) );
  OAI21X1 U583 ( .A(n4657), .B(n4744), .C(n2557), .Y(n1600) );
  OAI21X1 U586 ( .A(n4664), .B(n4742), .C(n3066), .Y(n1601) );
  OAI21X1 U588 ( .A(n4663), .B(n4742), .C(n3124), .Y(n1602) );
  OAI21X1 U590 ( .A(n4662), .B(n4742), .C(n3181), .Y(n1603) );
  OAI21X1 U592 ( .A(n4661), .B(n4742), .C(n3239), .Y(n1604) );
  OAI21X1 U594 ( .A(n4660), .B(n4742), .C(n3307), .Y(n1605) );
  OAI21X1 U596 ( .A(n4690), .B(n4742), .C(n3373), .Y(n1606) );
  OAI21X1 U598 ( .A(n4689), .B(n4742), .C(n3438), .Y(n1607) );
  OAI21X1 U600 ( .A(n4688), .B(n4742), .C(n3505), .Y(n1608) );
  OAI21X1 U602 ( .A(n4687), .B(n4742), .C(n2640), .Y(n1609) );
  OAI21X1 U604 ( .A(n4686), .B(n4742), .C(n3065), .Y(n1610) );
  OAI21X1 U606 ( .A(n4685), .B(n4742), .C(n2692), .Y(n1611) );
  OAI21X1 U608 ( .A(n4684), .B(n4742), .C(n2744), .Y(n1612) );
  OAI21X1 U610 ( .A(n4683), .B(n4742), .C(n2796), .Y(n1613) );
  OAI21X1 U612 ( .A(n4682), .B(n4742), .C(n3123), .Y(n1614) );
  OAI21X1 U614 ( .A(n4681), .B(n4743), .C(n3180), .Y(n1615) );
  OAI21X1 U616 ( .A(n4680), .B(n4742), .C(n3238), .Y(n1616) );
  OAI21X1 U618 ( .A(n4679), .B(n4743), .C(n3306), .Y(n1617) );
  OAI21X1 U620 ( .A(n4678), .B(n4742), .C(n3372), .Y(n1618) );
  OAI21X1 U622 ( .A(n4677), .B(n4743), .C(n3437), .Y(n1619) );
  OAI21X1 U624 ( .A(n4676), .B(n4742), .C(n3504), .Y(n1620) );
  OAI21X1 U626 ( .A(n4675), .B(n4743), .C(n2639), .Y(n1621) );
  OAI21X1 U628 ( .A(n4674), .B(n4742), .C(n2691), .Y(n1622) );
  OAI21X1 U630 ( .A(n4673), .B(n4743), .C(n2743), .Y(n1623) );
  OAI21X1 U632 ( .A(n4672), .B(n4742), .C(n2849), .Y(n1624) );
  OAI21X1 U634 ( .A(n4671), .B(n4742), .C(n2903), .Y(n1625) );
  OAI21X1 U636 ( .A(n4670), .B(n4742), .C(n2957), .Y(n1626) );
  OAI21X1 U638 ( .A(n4669), .B(n4742), .C(n3011), .Y(n1627) );
  OAI21X1 U640 ( .A(n4668), .B(n4742), .C(n2556), .Y(n1628) );
  OAI21X1 U642 ( .A(n4667), .B(n4742), .C(n2555), .Y(n1629) );
  OAI21X1 U644 ( .A(n4666), .B(n4743), .C(n2795), .Y(n1630) );
  OAI21X1 U646 ( .A(n4665), .B(n4742), .C(n2554), .Y(n1631) );
  OAI21X1 U648 ( .A(n4659), .B(n4742), .C(n2553), .Y(n1632) );
  OAI21X1 U650 ( .A(n4658), .B(n4742), .C(n2552), .Y(n1633) );
  OAI21X1 U652 ( .A(n4657), .B(n4742), .C(n2551), .Y(n1634) );
  NOR3X1 U655 ( .A(wr_ptr[3]), .B(wr_ptr[4]), .C(n1288), .Y(n190) );
  OAI21X1 U656 ( .A(n4664), .B(n4740), .C(n3010), .Y(n1635) );
  OAI21X1 U658 ( .A(n4663), .B(n4741), .C(n2956), .Y(n1636) );
  OAI21X1 U660 ( .A(n4662), .B(n4740), .C(n2902), .Y(n1637) );
  OAI21X1 U662 ( .A(n4661), .B(n4741), .C(n2848), .Y(n1638) );
  OAI21X1 U664 ( .A(n4660), .B(n4740), .C(n2794), .Y(n1639) );
  OAI21X1 U666 ( .A(n4690), .B(n4741), .C(n2742), .Y(n1640) );
  OAI21X1 U668 ( .A(n4689), .B(n4740), .C(n2690), .Y(n1641) );
  OAI21X1 U670 ( .A(n4688), .B(n4741), .C(n2638), .Y(n1642) );
  OAI21X1 U672 ( .A(n4687), .B(n4740), .C(n3503), .Y(n1643) );
  OAI21X1 U674 ( .A(n4686), .B(n4741), .C(n3009), .Y(n1644) );
  OAI21X1 U676 ( .A(n4685), .B(n4740), .C(n3436), .Y(n1645) );
  OAI21X1 U678 ( .A(n4684), .B(n4741), .C(n3371), .Y(n1646) );
  OAI21X1 U680 ( .A(n4683), .B(n4740), .C(n3305), .Y(n1647) );
  OAI21X1 U682 ( .A(n4682), .B(n4740), .C(n2955), .Y(n1648) );
  OAI21X1 U684 ( .A(n4681), .B(n4741), .C(n2901), .Y(n1649) );
  OAI21X1 U686 ( .A(n4680), .B(n4741), .C(n2847), .Y(n1650) );
  OAI21X1 U688 ( .A(n4679), .B(n4740), .C(n2793), .Y(n1651) );
  OAI21X1 U690 ( .A(n4678), .B(n4741), .C(n2741), .Y(n1652) );
  OAI21X1 U692 ( .A(n4677), .B(n4740), .C(n2689), .Y(n1653) );
  OAI21X1 U694 ( .A(n4676), .B(n4741), .C(n2637), .Y(n1654) );
  OAI21X1 U696 ( .A(n4675), .B(n4740), .C(n3502), .Y(n1655) );
  OAI21X1 U698 ( .A(n4674), .B(n4740), .C(n3435), .Y(n1656) );
  OAI21X1 U700 ( .A(n4673), .B(n4740), .C(n3370), .Y(n1657) );
  OAI21X1 U702 ( .A(n4672), .B(n4740), .C(n3237), .Y(n1658) );
  OAI21X1 U704 ( .A(n4671), .B(n4740), .C(n3179), .Y(n1659) );
  OAI21X1 U706 ( .A(n4670), .B(n4740), .C(n3122), .Y(n1660) );
  OAI21X1 U708 ( .A(n4669), .B(n4740), .C(n3064), .Y(n1661) );
  OAI21X1 U710 ( .A(n4668), .B(n4740), .C(n2550), .Y(n1662) );
  OAI21X1 U712 ( .A(n4667), .B(n4740), .C(n2549), .Y(n1663) );
  OAI21X1 U714 ( .A(n4666), .B(n4740), .C(n3304), .Y(n1664) );
  OAI21X1 U716 ( .A(n4665), .B(n4740), .C(n2548), .Y(n1665) );
  OAI21X1 U718 ( .A(n4659), .B(n4740), .C(n2547), .Y(n1666) );
  OAI21X1 U720 ( .A(n4658), .B(n4740), .C(n2546), .Y(n1667) );
  OAI21X1 U722 ( .A(n4657), .B(n4740), .C(n2545), .Y(n1668) );
  OAI21X1 U725 ( .A(n4664), .B(n4738), .C(n2954), .Y(n1669) );
  OAI21X1 U727 ( .A(n4663), .B(n4739), .C(n3008), .Y(n1670) );
  OAI21X1 U729 ( .A(n4662), .B(n4738), .C(n2846), .Y(n1671) );
  OAI21X1 U731 ( .A(n4661), .B(n4739), .C(n2900), .Y(n1672) );
  OAI21X1 U733 ( .A(n4660), .B(n4738), .C(n2740), .Y(n1673) );
  OAI21X1 U735 ( .A(n4690), .B(n4739), .C(n2792), .Y(n1674) );
  OAI21X1 U737 ( .A(n4689), .B(n4738), .C(n2636), .Y(n1675) );
  OAI21X1 U739 ( .A(n4688), .B(n4739), .C(n2688), .Y(n1676) );
  OAI21X1 U741 ( .A(n4687), .B(n4738), .C(n3434), .Y(n1677) );
  OAI21X1 U743 ( .A(n4686), .B(n4739), .C(n2953), .Y(n1678) );
  OAI21X1 U745 ( .A(n4685), .B(n4738), .C(n3501), .Y(n1679) );
  OAI21X1 U747 ( .A(n4684), .B(n4739), .C(n3303), .Y(n1680) );
  OAI21X1 U749 ( .A(n4683), .B(n4738), .C(n3369), .Y(n1681) );
  OAI21X1 U751 ( .A(n4682), .B(n4738), .C(n3007), .Y(n1682) );
  OAI21X1 U753 ( .A(n4681), .B(n4739), .C(n2845), .Y(n1683) );
  OAI21X1 U755 ( .A(n4680), .B(n4739), .C(n2899), .Y(n1684) );
  OAI21X1 U757 ( .A(n4679), .B(n4738), .C(n2739), .Y(n1685) );
  OAI21X1 U759 ( .A(n4678), .B(n4739), .C(n2791), .Y(n1686) );
  OAI21X1 U761 ( .A(n4677), .B(n4738), .C(n2635), .Y(n1687) );
  OAI21X1 U763 ( .A(n4676), .B(n4739), .C(n2687), .Y(n1688) );
  OAI21X1 U765 ( .A(n4675), .B(n4738), .C(n3433), .Y(n1689) );
  OAI21X1 U767 ( .A(n4674), .B(n4738), .C(n3500), .Y(n1690) );
  OAI21X1 U769 ( .A(n4673), .B(n4738), .C(n3302), .Y(n1691) );
  OAI21X1 U771 ( .A(n4672), .B(n4738), .C(n3178), .Y(n1692) );
  OAI21X1 U773 ( .A(n4671), .B(n4738), .C(n3236), .Y(n1693) );
  OAI21X1 U775 ( .A(n4670), .B(n4738), .C(n3063), .Y(n1694) );
  OAI21X1 U777 ( .A(n4669), .B(n4738), .C(n3121), .Y(n1695) );
  OAI21X1 U779 ( .A(n4668), .B(n4738), .C(n2544), .Y(n1696) );
  OAI21X1 U781 ( .A(n4667), .B(n4738), .C(n2543), .Y(n1697) );
  OAI21X1 U783 ( .A(n4666), .B(n4738), .C(n3368), .Y(n1698) );
  OAI21X1 U785 ( .A(n4665), .B(n4738), .C(n2542), .Y(n1699) );
  OAI21X1 U787 ( .A(n4659), .B(n4738), .C(n2541), .Y(n1700) );
  OAI21X1 U789 ( .A(n4658), .B(n4738), .C(n2540), .Y(n1701) );
  OAI21X1 U791 ( .A(n4657), .B(n4738), .C(n2539), .Y(n1702) );
  OAI21X1 U794 ( .A(n4664), .B(n4736), .C(n2898), .Y(n1703) );
  OAI21X1 U796 ( .A(n4663), .B(n4737), .C(n2844), .Y(n1704) );
  OAI21X1 U798 ( .A(n4662), .B(n4736), .C(n3006), .Y(n1705) );
  OAI21X1 U800 ( .A(n4661), .B(n4737), .C(n2952), .Y(n1706) );
  OAI21X1 U802 ( .A(n4660), .B(n4736), .C(n2686), .Y(n1707) );
  OAI21X1 U804 ( .A(n4690), .B(n4737), .C(n2634), .Y(n1708) );
  OAI21X1 U806 ( .A(n4689), .B(n4736), .C(n2790), .Y(n1709) );
  OAI21X1 U808 ( .A(n4688), .B(n4737), .C(n2738), .Y(n1710) );
  OAI21X1 U810 ( .A(n4687), .B(n4736), .C(n3367), .Y(n1711) );
  OAI21X1 U812 ( .A(n4686), .B(n4737), .C(n2897), .Y(n1712) );
  OAI21X1 U814 ( .A(n4685), .B(n4736), .C(n3301), .Y(n1713) );
  OAI21X1 U816 ( .A(n4684), .B(n4737), .C(n3499), .Y(n1714) );
  OAI21X1 U818 ( .A(n4683), .B(n4736), .C(n3432), .Y(n1715) );
  OAI21X1 U820 ( .A(n4682), .B(n4736), .C(n2843), .Y(n1716) );
  OAI21X1 U822 ( .A(n4681), .B(n4737), .C(n3005), .Y(n1717) );
  OAI21X1 U824 ( .A(n4680), .B(n4737), .C(n2951), .Y(n1718) );
  OAI21X1 U826 ( .A(n4679), .B(n4736), .C(n2685), .Y(n1719) );
  OAI21X1 U828 ( .A(n4678), .B(n4737), .C(n2633), .Y(n1720) );
  OAI21X1 U830 ( .A(n4677), .B(n4736), .C(n2789), .Y(n1721) );
  OAI21X1 U832 ( .A(n4676), .B(n4737), .C(n2737), .Y(n1722) );
  OAI21X1 U834 ( .A(n4675), .B(n4736), .C(n3366), .Y(n1723) );
  OAI21X1 U836 ( .A(n4674), .B(n4736), .C(n3300), .Y(n1724) );
  OAI21X1 U838 ( .A(n4673), .B(n4736), .C(n3498), .Y(n1725) );
  OAI21X1 U840 ( .A(n4672), .B(n4736), .C(n3120), .Y(n1726) );
  OAI21X1 U842 ( .A(n4671), .B(n4736), .C(n3062), .Y(n1727) );
  OAI21X1 U844 ( .A(n4670), .B(n4736), .C(n3235), .Y(n1728) );
  OAI21X1 U846 ( .A(n4669), .B(n4736), .C(n3177), .Y(n1729) );
  OAI21X1 U848 ( .A(n4668), .B(n4736), .C(n2538), .Y(n1730) );
  OAI21X1 U850 ( .A(n4667), .B(n4736), .C(n2537), .Y(n1731) );
  OAI21X1 U852 ( .A(n4666), .B(n4736), .C(n3431), .Y(n1732) );
  OAI21X1 U854 ( .A(n4665), .B(n4736), .C(n2536), .Y(n1733) );
  OAI21X1 U856 ( .A(n4659), .B(n4736), .C(n2535), .Y(n1734) );
  OAI21X1 U858 ( .A(n4658), .B(n4736), .C(n2534), .Y(n1735) );
  OAI21X1 U860 ( .A(n4657), .B(n4736), .C(n2533), .Y(n1736) );
  OAI21X1 U863 ( .A(n4664), .B(n4734), .C(n2842), .Y(n1737) );
  OAI21X1 U865 ( .A(n4663), .B(n4735), .C(n2896), .Y(n1738) );
  OAI21X1 U867 ( .A(n4662), .B(n4734), .C(n2950), .Y(n1739) );
  OAI21X1 U869 ( .A(n4661), .B(n4735), .C(n3004), .Y(n1740) );
  OAI21X1 U871 ( .A(n4660), .B(n4734), .C(n2632), .Y(n1741) );
  OAI21X1 U873 ( .A(n4690), .B(n4735), .C(n2684), .Y(n1742) );
  OAI21X1 U875 ( .A(n4689), .B(n4734), .C(n2736), .Y(n1743) );
  OAI21X1 U877 ( .A(n4688), .B(n4735), .C(n2788), .Y(n1744) );
  OAI21X1 U879 ( .A(n4687), .B(n4734), .C(n3299), .Y(n1745) );
  OAI21X1 U881 ( .A(n4686), .B(n4735), .C(n2841), .Y(n1746) );
  OAI21X1 U883 ( .A(n4685), .B(n4734), .C(n3365), .Y(n1747) );
  OAI21X1 U885 ( .A(n4684), .B(n4735), .C(n3430), .Y(n1748) );
  OAI21X1 U887 ( .A(n4683), .B(n4734), .C(n3497), .Y(n1749) );
  OAI21X1 U889 ( .A(n4682), .B(n4734), .C(n2895), .Y(n1750) );
  OAI21X1 U891 ( .A(n4681), .B(n4735), .C(n2949), .Y(n1751) );
  OAI21X1 U893 ( .A(n4680), .B(n4735), .C(n3003), .Y(n1752) );
  OAI21X1 U895 ( .A(n4679), .B(n4734), .C(n2631), .Y(n1753) );
  OAI21X1 U897 ( .A(n4678), .B(n4735), .C(n2683), .Y(n1754) );
  OAI21X1 U899 ( .A(n4677), .B(n4734), .C(n2735), .Y(n1755) );
  OAI21X1 U901 ( .A(n4676), .B(n4735), .C(n2787), .Y(n1756) );
  OAI21X1 U903 ( .A(n4675), .B(n4734), .C(n3298), .Y(n1757) );
  OAI21X1 U905 ( .A(n4674), .B(n4734), .C(n3364), .Y(n1758) );
  OAI21X1 U907 ( .A(n4673), .B(n4734), .C(n3429), .Y(n1759) );
  OAI21X1 U909 ( .A(n4672), .B(n4734), .C(n3061), .Y(n1760) );
  OAI21X1 U911 ( .A(n4671), .B(n4734), .C(n3119), .Y(n1761) );
  OAI21X1 U913 ( .A(n4670), .B(n4734), .C(n3176), .Y(n1762) );
  OAI21X1 U915 ( .A(n4669), .B(n4734), .C(n3234), .Y(n1763) );
  OAI21X1 U917 ( .A(n4668), .B(n4734), .C(n2532), .Y(n1764) );
  OAI21X1 U919 ( .A(n4667), .B(n4734), .C(n2531), .Y(n1765) );
  OAI21X1 U921 ( .A(n4666), .B(n4734), .C(n3496), .Y(n1766) );
  OAI21X1 U923 ( .A(n4665), .B(n4734), .C(n2530), .Y(n1767) );
  OAI21X1 U925 ( .A(n4659), .B(n4734), .C(n2529), .Y(n1768) );
  OAI21X1 U927 ( .A(n4658), .B(n4734), .C(n2528), .Y(n1769) );
  OAI21X1 U929 ( .A(n4657), .B(n4734), .C(n2527), .Y(n1770) );
  OAI21X1 U932 ( .A(n4664), .B(n4732), .C(n2786), .Y(n1771) );
  OAI21X1 U934 ( .A(n4663), .B(n4733), .C(n2734), .Y(n1772) );
  OAI21X1 U936 ( .A(n4662), .B(n4732), .C(n2682), .Y(n1773) );
  OAI21X1 U938 ( .A(n4661), .B(n4733), .C(n2630), .Y(n1774) );
  OAI21X1 U940 ( .A(n4660), .B(n4732), .C(n3002), .Y(n1775) );
  OAI21X1 U942 ( .A(n4690), .B(n4733), .C(n2948), .Y(n1776) );
  OAI21X1 U944 ( .A(n4689), .B(n4732), .C(n2894), .Y(n1777) );
  OAI21X1 U946 ( .A(n4688), .B(n4733), .C(n2840), .Y(n1778) );
  OAI21X1 U948 ( .A(n4687), .B(n4732), .C(n3233), .Y(n1779) );
  OAI21X1 U950 ( .A(n4686), .B(n4733), .C(n2785), .Y(n1780) );
  OAI21X1 U952 ( .A(n4685), .B(n4732), .C(n3175), .Y(n1781) );
  OAI21X1 U954 ( .A(n4684), .B(n4733), .C(n3118), .Y(n1782) );
  OAI21X1 U956 ( .A(n4683), .B(n4732), .C(n3060), .Y(n1783) );
  OAI21X1 U958 ( .A(n4682), .B(n4732), .C(n2733), .Y(n1784) );
  OAI21X1 U960 ( .A(n4681), .B(n4733), .C(n2681), .Y(n1785) );
  OAI21X1 U962 ( .A(n4680), .B(n4733), .C(n2629), .Y(n1786) );
  OAI21X1 U964 ( .A(n4679), .B(n4732), .C(n3001), .Y(n1787) );
  OAI21X1 U966 ( .A(n4678), .B(n4733), .C(n2947), .Y(n1788) );
  OAI21X1 U968 ( .A(n4677), .B(n4732), .C(n2893), .Y(n1789) );
  OAI21X1 U970 ( .A(n4676), .B(n4733), .C(n2839), .Y(n1790) );
  OAI21X1 U972 ( .A(n4675), .B(n4732), .C(n3232), .Y(n1791) );
  OAI21X1 U974 ( .A(n4674), .B(n4732), .C(n3174), .Y(n1792) );
  OAI21X1 U976 ( .A(n4673), .B(n4732), .C(n3117), .Y(n1793) );
  OAI21X1 U978 ( .A(n4672), .B(n4732), .C(n3495), .Y(n1794) );
  OAI21X1 U980 ( .A(n4671), .B(n4732), .C(n3428), .Y(n1795) );
  OAI21X1 U982 ( .A(n4670), .B(n4732), .C(n3363), .Y(n1796) );
  OAI21X1 U984 ( .A(n4669), .B(n4732), .C(n3297), .Y(n1797) );
  OAI21X1 U986 ( .A(n4668), .B(n4732), .C(n2526), .Y(n1798) );
  OAI21X1 U988 ( .A(n4667), .B(n4732), .C(n2525), .Y(n1799) );
  OAI21X1 U990 ( .A(n4666), .B(n4732), .C(n3059), .Y(n1800) );
  OAI21X1 U992 ( .A(n4665), .B(n4732), .C(n2524), .Y(n1801) );
  OAI21X1 U994 ( .A(n4659), .B(n4732), .C(n2523), .Y(n1802) );
  OAI21X1 U996 ( .A(n4658), .B(n4732), .C(n2522), .Y(n1803) );
  OAI21X1 U998 ( .A(n4657), .B(n4732), .C(n2521), .Y(n1804) );
  OAI21X1 U1001 ( .A(n4664), .B(n4730), .C(n3494), .Y(n1805) );
  OAI21X1 U1003 ( .A(n4663), .B(n4731), .C(n3427), .Y(n1806) );
  OAI21X1 U1005 ( .A(n4662), .B(n4730), .C(n3362), .Y(n1807) );
  OAI21X1 U1007 ( .A(n4661), .B(n4731), .C(n3296), .Y(n1808) );
  OAI21X1 U1009 ( .A(n4660), .B(n4730), .C(n3231), .Y(n1809) );
  OAI21X1 U1011 ( .A(n4690), .B(n4731), .C(n3173), .Y(n1810) );
  OAI21X1 U1013 ( .A(n4689), .B(n4730), .C(n3116), .Y(n1811) );
  OAI21X1 U1015 ( .A(n4688), .B(n4731), .C(n3058), .Y(n1812) );
  OAI21X1 U1017 ( .A(n4687), .B(n4730), .C(n3000), .Y(n1813) );
  OAI21X1 U1019 ( .A(n4686), .B(n4731), .C(n3493), .Y(n1814) );
  OAI21X1 U1021 ( .A(n4685), .B(n4730), .C(n2946), .Y(n1815) );
  OAI21X1 U1023 ( .A(n4684), .B(n4731), .C(n2892), .Y(n1816) );
  OAI21X1 U1025 ( .A(n4683), .B(n4730), .C(n2838), .Y(n1817) );
  OAI21X1 U1027 ( .A(n4682), .B(n4730), .C(n3426), .Y(n1818) );
  OAI21X1 U1029 ( .A(n4681), .B(n4731), .C(n3361), .Y(n1819) );
  OAI21X1 U1031 ( .A(n4680), .B(n4731), .C(n3295), .Y(n1820) );
  OAI21X1 U1033 ( .A(n4679), .B(n4730), .C(n3230), .Y(n1821) );
  OAI21X1 U1035 ( .A(n4678), .B(n4731), .C(n3172), .Y(n1822) );
  OAI21X1 U1037 ( .A(n4677), .B(n4730), .C(n3115), .Y(n1823) );
  OAI21X1 U1039 ( .A(n4676), .B(n4731), .C(n3057), .Y(n1824) );
  OAI21X1 U1041 ( .A(n4675), .B(n4730), .C(n2999), .Y(n1825) );
  OAI21X1 U1043 ( .A(n4674), .B(n4730), .C(n2945), .Y(n1826) );
  OAI21X1 U1045 ( .A(n4673), .B(n4730), .C(n2891), .Y(n1827) );
  OAI21X1 U1047 ( .A(n4672), .B(n4730), .C(n2784), .Y(n1828) );
  OAI21X1 U1049 ( .A(n4671), .B(n4730), .C(n2732), .Y(n1829) );
  OAI21X1 U1051 ( .A(n4670), .B(n4730), .C(n2680), .Y(n1830) );
  OAI21X1 U1053 ( .A(n4669), .B(n4730), .C(n2628), .Y(n1831) );
  OAI21X1 U1055 ( .A(n4668), .B(n4730), .C(n2520), .Y(n1832) );
  OAI21X1 U1057 ( .A(n4667), .B(n4730), .C(n2519), .Y(n1833) );
  OAI21X1 U1059 ( .A(n4666), .B(n4730), .C(n2837), .Y(n1834) );
  OAI21X1 U1061 ( .A(n4665), .B(n4730), .C(n2518), .Y(n1835) );
  OAI21X1 U1063 ( .A(n4659), .B(n4730), .C(n2517), .Y(n1836) );
  OAI21X1 U1065 ( .A(n4658), .B(n4730), .C(n2516), .Y(n1837) );
  OAI21X1 U1067 ( .A(n4657), .B(n4730), .C(n2515), .Y(n1838) );
  OAI21X1 U1070 ( .A(n4664), .B(n4728), .C(n3425), .Y(n1839) );
  OAI21X1 U1072 ( .A(n4663), .B(n4729), .C(n3492), .Y(n1840) );
  OAI21X1 U1074 ( .A(n4662), .B(n4728), .C(n3294), .Y(n1841) );
  OAI21X1 U1076 ( .A(n4661), .B(n4729), .C(n3360), .Y(n1842) );
  OAI21X1 U1078 ( .A(n4660), .B(n4728), .C(n3171), .Y(n1843) );
  OAI21X1 U1080 ( .A(n4690), .B(n4729), .C(n3229), .Y(n1844) );
  OAI21X1 U1082 ( .A(n4689), .B(n4728), .C(n3056), .Y(n1845) );
  OAI21X1 U1084 ( .A(n4688), .B(n4729), .C(n3114), .Y(n1846) );
  OAI21X1 U1086 ( .A(n4687), .B(n4728), .C(n2944), .Y(n1847) );
  OAI21X1 U1088 ( .A(n4686), .B(n4729), .C(n3424), .Y(n1848) );
  OAI21X1 U1090 ( .A(n4685), .B(n4728), .C(n2998), .Y(n1849) );
  OAI21X1 U1092 ( .A(n4684), .B(n4729), .C(n2836), .Y(n1850) );
  OAI21X1 U1094 ( .A(n4683), .B(n4728), .C(n2890), .Y(n1851) );
  OAI21X1 U1096 ( .A(n4682), .B(n4728), .C(n3491), .Y(n1852) );
  OAI21X1 U1098 ( .A(n4681), .B(n4729), .C(n3293), .Y(n1853) );
  OAI21X1 U1100 ( .A(n4680), .B(n4729), .C(n3359), .Y(n1854) );
  OAI21X1 U1102 ( .A(n4679), .B(n4728), .C(n3170), .Y(n1855) );
  OAI21X1 U1104 ( .A(n4678), .B(n4729), .C(n3228), .Y(n1856) );
  OAI21X1 U1106 ( .A(n4677), .B(n4728), .C(n3055), .Y(n1857) );
  OAI21X1 U1108 ( .A(n4676), .B(n4729), .C(n3113), .Y(n1858) );
  OAI21X1 U1110 ( .A(n4675), .B(n4728), .C(n2943), .Y(n1859) );
  OAI21X1 U1112 ( .A(n4674), .B(n4728), .C(n2997), .Y(n1860) );
  OAI21X1 U1114 ( .A(n4673), .B(n4728), .C(n2835), .Y(n1861) );
  OAI21X1 U1116 ( .A(n4672), .B(n4728), .C(n2731), .Y(n1862) );
  OAI21X1 U1118 ( .A(n4671), .B(n4728), .C(n2783), .Y(n1863) );
  OAI21X1 U1120 ( .A(n4670), .B(n4728), .C(n2627), .Y(n1864) );
  OAI21X1 U1122 ( .A(n4669), .B(n4728), .C(n2679), .Y(n1865) );
  OAI21X1 U1124 ( .A(n4668), .B(n4728), .C(n2514), .Y(n1866) );
  OAI21X1 U1126 ( .A(n4667), .B(n4728), .C(n2513), .Y(n1867) );
  OAI21X1 U1128 ( .A(n4666), .B(n4728), .C(n2889), .Y(n1868) );
  OAI21X1 U1130 ( .A(n4665), .B(n4728), .C(n2512), .Y(n1869) );
  OAI21X1 U1132 ( .A(n4659), .B(n4728), .C(n2511), .Y(n1870) );
  OAI21X1 U1134 ( .A(n4658), .B(n4728), .C(n2510), .Y(n1871) );
  OAI21X1 U1136 ( .A(n4657), .B(n4728), .C(n2509), .Y(n1872) );
  OAI21X1 U1139 ( .A(n4664), .B(n4726), .C(n3358), .Y(n1873) );
  OAI21X1 U1141 ( .A(n4663), .B(n4727), .C(n3292), .Y(n1874) );
  OAI21X1 U1143 ( .A(n4662), .B(n4726), .C(n3490), .Y(n1875) );
  OAI21X1 U1145 ( .A(n4661), .B(n4727), .C(n3423), .Y(n1876) );
  OAI21X1 U1147 ( .A(n4660), .B(n4726), .C(n3112), .Y(n1877) );
  OAI21X1 U1149 ( .A(n4690), .B(n4727), .C(n3054), .Y(n1878) );
  OAI21X1 U1151 ( .A(n4689), .B(n4726), .C(n3227), .Y(n1879) );
  OAI21X1 U1153 ( .A(n4688), .B(n4727), .C(n3169), .Y(n1880) );
  OAI21X1 U1155 ( .A(n4687), .B(n4726), .C(n2888), .Y(n1881) );
  OAI21X1 U1157 ( .A(n4686), .B(n4727), .C(n3357), .Y(n1882) );
  OAI21X1 U1159 ( .A(n4685), .B(n4726), .C(n2834), .Y(n1883) );
  OAI21X1 U1161 ( .A(n4684), .B(n4727), .C(n2996), .Y(n1884) );
  OAI21X1 U1163 ( .A(n4683), .B(n4726), .C(n2942), .Y(n1885) );
  OAI21X1 U1165 ( .A(n4682), .B(n4726), .C(n3291), .Y(n1886) );
  OAI21X1 U1167 ( .A(n4681), .B(n4727), .C(n3489), .Y(n1887) );
  OAI21X1 U1169 ( .A(n4680), .B(n4727), .C(n3422), .Y(n1888) );
  OAI21X1 U1171 ( .A(n4679), .B(n4726), .C(n3111), .Y(n1889) );
  OAI21X1 U1173 ( .A(n4678), .B(n4727), .C(n3053), .Y(n1890) );
  OAI21X1 U1175 ( .A(n4677), .B(n4726), .C(n3226), .Y(n1891) );
  OAI21X1 U1177 ( .A(n4676), .B(n4727), .C(n3168), .Y(n1892) );
  OAI21X1 U1179 ( .A(n4675), .B(n4726), .C(n2887), .Y(n1893) );
  OAI21X1 U1181 ( .A(n4674), .B(n4726), .C(n2833), .Y(n1894) );
  OAI21X1 U1183 ( .A(n4673), .B(n4726), .C(n2995), .Y(n1895) );
  OAI21X1 U1185 ( .A(n4672), .B(n4726), .C(n2678), .Y(n1896) );
  OAI21X1 U1187 ( .A(n4671), .B(n4726), .C(n2626), .Y(n1897) );
  OAI21X1 U1189 ( .A(n4670), .B(n4726), .C(n2782), .Y(n1898) );
  OAI21X1 U1191 ( .A(n4669), .B(n4726), .C(n2730), .Y(n1899) );
  OAI21X1 U1193 ( .A(n4668), .B(n4726), .C(n2508), .Y(n1900) );
  OAI21X1 U1195 ( .A(n4667), .B(n4726), .C(n2507), .Y(n1901) );
  OAI21X1 U1197 ( .A(n4666), .B(n4726), .C(n2941), .Y(n1902) );
  OAI21X1 U1199 ( .A(n4665), .B(n4726), .C(n2506), .Y(n1903) );
  OAI21X1 U1201 ( .A(n4659), .B(n4726), .C(n2505), .Y(n1904) );
  OAI21X1 U1203 ( .A(n4658), .B(n4726), .C(n2504), .Y(n1905) );
  OAI21X1 U1205 ( .A(n4657), .B(n4726), .C(n2503), .Y(n1906) );
  NOR3X1 U1208 ( .A(n1288), .B(wr_ptr[4]), .C(n4811), .Y(n478) );
  OAI21X1 U1209 ( .A(n4664), .B(n4724), .C(n3290), .Y(n1907) );
  OAI21X1 U1211 ( .A(n4663), .B(n4725), .C(n3356), .Y(n1908) );
  OAI21X1 U1213 ( .A(n4662), .B(n4724), .C(n3421), .Y(n1909) );
  OAI21X1 U1215 ( .A(n4661), .B(n4725), .C(n3488), .Y(n1910) );
  OAI21X1 U1217 ( .A(n4660), .B(n4724), .C(n3052), .Y(n1911) );
  OAI21X1 U1219 ( .A(n4690), .B(n4725), .C(n3110), .Y(n1912) );
  OAI21X1 U1221 ( .A(n4689), .B(n4724), .C(n3167), .Y(n1913) );
  OAI21X1 U1223 ( .A(n4688), .B(n4725), .C(n3225), .Y(n1914) );
  OAI21X1 U1225 ( .A(n4687), .B(n4724), .C(n2832), .Y(n1915) );
  OAI21X1 U1227 ( .A(n4686), .B(n4725), .C(n3289), .Y(n1916) );
  OAI21X1 U1229 ( .A(n4685), .B(n4724), .C(n2886), .Y(n1917) );
  OAI21X1 U1231 ( .A(n4684), .B(n4725), .C(n2940), .Y(n1918) );
  OAI21X1 U1233 ( .A(n4683), .B(n4724), .C(n2994), .Y(n1919) );
  OAI21X1 U1235 ( .A(n4682), .B(n4724), .C(n3355), .Y(n1920) );
  OAI21X1 U1237 ( .A(n4681), .B(n4725), .C(n3420), .Y(n1921) );
  OAI21X1 U1239 ( .A(n4680), .B(n4725), .C(n3487), .Y(n1922) );
  OAI21X1 U1241 ( .A(n4679), .B(n4724), .C(n3051), .Y(n1923) );
  OAI21X1 U1243 ( .A(n4678), .B(n4725), .C(n3109), .Y(n1924) );
  OAI21X1 U1245 ( .A(n4677), .B(n4724), .C(n3166), .Y(n1925) );
  OAI21X1 U1247 ( .A(n4676), .B(n4725), .C(n3224), .Y(n1926) );
  OAI21X1 U1249 ( .A(n4675), .B(n4724), .C(n2831), .Y(n1927) );
  OAI21X1 U1251 ( .A(n4674), .B(n4724), .C(n2885), .Y(n1928) );
  OAI21X1 U1253 ( .A(n4673), .B(n4724), .C(n2939), .Y(n1929) );
  OAI21X1 U1255 ( .A(n4672), .B(n4724), .C(n2625), .Y(n1930) );
  OAI21X1 U1257 ( .A(n4671), .B(n4724), .C(n2677), .Y(n1931) );
  OAI21X1 U1259 ( .A(n4670), .B(n4724), .C(n2729), .Y(n1932) );
  OAI21X1 U1261 ( .A(n4669), .B(n4724), .C(n2781), .Y(n1933) );
  OAI21X1 U1263 ( .A(n4668), .B(n4724), .C(n2502), .Y(n1934) );
  OAI21X1 U1265 ( .A(n4667), .B(n4724), .C(n2501), .Y(n1935) );
  OAI21X1 U1267 ( .A(n4666), .B(n4724), .C(n2993), .Y(n1936) );
  OAI21X1 U1269 ( .A(n4665), .B(n4724), .C(n2500), .Y(n1937) );
  OAI21X1 U1271 ( .A(n4659), .B(n4724), .C(n2499), .Y(n1938) );
  OAI21X1 U1273 ( .A(n4658), .B(n4724), .C(n2498), .Y(n1939) );
  OAI21X1 U1275 ( .A(n4657), .B(n4724), .C(n2497), .Y(n1940) );
  OAI21X1 U1278 ( .A(n4664), .B(n4722), .C(n3223), .Y(n1941) );
  OAI21X1 U1280 ( .A(n4663), .B(n4723), .C(n3165), .Y(n1942) );
  OAI21X1 U1282 ( .A(n4662), .B(n4722), .C(n3108), .Y(n1943) );
  OAI21X1 U1284 ( .A(n4661), .B(n4723), .C(n3050), .Y(n1944) );
  OAI21X1 U1286 ( .A(n4660), .B(n4722), .C(n3486), .Y(n1945) );
  OAI21X1 U1288 ( .A(n4690), .B(n4723), .C(n3419), .Y(n1946) );
  OAI21X1 U1290 ( .A(n4689), .B(n4722), .C(n3354), .Y(n1947) );
  OAI21X1 U1292 ( .A(n4688), .B(n4723), .C(n3288), .Y(n1948) );
  OAI21X1 U1294 ( .A(n4687), .B(n4722), .C(n2780), .Y(n1949) );
  OAI21X1 U1296 ( .A(n4686), .B(n4723), .C(n3222), .Y(n1950) );
  OAI21X1 U1298 ( .A(n4685), .B(n4722), .C(n2728), .Y(n1951) );
  OAI21X1 U1300 ( .A(n4684), .B(n4723), .C(n2676), .Y(n1952) );
  OAI21X1 U1302 ( .A(n4683), .B(n4722), .C(n2624), .Y(n1953) );
  OAI21X1 U1304 ( .A(n4682), .B(n4722), .C(n3164), .Y(n1954) );
  OAI21X1 U1306 ( .A(n4681), .B(n4723), .C(n3107), .Y(n1955) );
  OAI21X1 U1308 ( .A(n4680), .B(n4723), .C(n3049), .Y(n1956) );
  OAI21X1 U1310 ( .A(n4679), .B(n4722), .C(n3485), .Y(n1957) );
  OAI21X1 U1312 ( .A(n4678), .B(n4723), .C(n3418), .Y(n1958) );
  OAI21X1 U1314 ( .A(n4677), .B(n4722), .C(n3353), .Y(n1959) );
  OAI21X1 U1316 ( .A(n4676), .B(n4723), .C(n3287), .Y(n1960) );
  OAI21X1 U1318 ( .A(n4675), .B(n4722), .C(n2779), .Y(n1961) );
  OAI21X1 U1320 ( .A(n4674), .B(n4722), .C(n2727), .Y(n1962) );
  OAI21X1 U1322 ( .A(n4673), .B(n4722), .C(n2675), .Y(n1963) );
  OAI21X1 U1324 ( .A(n4672), .B(n4722), .C(n2992), .Y(n1964) );
  OAI21X1 U1326 ( .A(n4671), .B(n4722), .C(n2938), .Y(n1965) );
  OAI21X1 U1328 ( .A(n4670), .B(n4722), .C(n2884), .Y(n1966) );
  OAI21X1 U1330 ( .A(n4669), .B(n4722), .C(n2830), .Y(n1967) );
  OAI21X1 U1332 ( .A(n4668), .B(n4722), .C(n2496), .Y(n1968) );
  OAI21X1 U1334 ( .A(n4667), .B(n4722), .C(n2495), .Y(n1969) );
  OAI21X1 U1336 ( .A(n4666), .B(n4722), .C(n2623), .Y(n1970) );
  OAI21X1 U1338 ( .A(n4665), .B(n4722), .C(n2494), .Y(n1971) );
  OAI21X1 U1340 ( .A(n4659), .B(n4722), .C(n2493), .Y(n1972) );
  OAI21X1 U1342 ( .A(n4658), .B(n4722), .C(n2492), .Y(n1973) );
  OAI21X1 U1344 ( .A(n4657), .B(n4722), .C(n2491), .Y(n1974) );
  OAI21X1 U1347 ( .A(n4664), .B(n4720), .C(n3163), .Y(n1975) );
  OAI21X1 U1349 ( .A(n4663), .B(n4721), .C(n3221), .Y(n1976) );
  OAI21X1 U1351 ( .A(n4662), .B(n4720), .C(n3048), .Y(n1977) );
  OAI21X1 U1353 ( .A(n4661), .B(n4721), .C(n3106), .Y(n1978) );
  OAI21X1 U1355 ( .A(n4660), .B(n4720), .C(n3417), .Y(n1979) );
  OAI21X1 U1357 ( .A(n4690), .B(n4721), .C(n3484), .Y(n1980) );
  OAI21X1 U1359 ( .A(n4689), .B(n4720), .C(n3286), .Y(n1981) );
  OAI21X1 U1361 ( .A(n4688), .B(n4721), .C(n3352), .Y(n1982) );
  OAI21X1 U1363 ( .A(n4687), .B(n4720), .C(n2726), .Y(n1983) );
  OAI21X1 U1365 ( .A(n4686), .B(n4721), .C(n3162), .Y(n1984) );
  OAI21X1 U1367 ( .A(n4685), .B(n4720), .C(n2778), .Y(n1985) );
  OAI21X1 U1369 ( .A(n4684), .B(n4721), .C(n2622), .Y(n1986) );
  OAI21X1 U1371 ( .A(n4683), .B(n4720), .C(n2674), .Y(n1987) );
  OAI21X1 U1373 ( .A(n4682), .B(n4720), .C(n3220), .Y(n1988) );
  OAI21X1 U1375 ( .A(n4681), .B(n4721), .C(n3047), .Y(n1989) );
  OAI21X1 U1377 ( .A(n4680), .B(n4721), .C(n3105), .Y(n1990) );
  OAI21X1 U1379 ( .A(n4679), .B(n4720), .C(n3416), .Y(n1991) );
  OAI21X1 U1381 ( .A(n4678), .B(n4721), .C(n3483), .Y(n1992) );
  OAI21X1 U1383 ( .A(n4677), .B(n4720), .C(n3285), .Y(n1993) );
  OAI21X1 U1385 ( .A(n4676), .B(n4721), .C(n3351), .Y(n1994) );
  OAI21X1 U1387 ( .A(n4675), .B(n4720), .C(n2725), .Y(n1995) );
  OAI21X1 U1389 ( .A(n4674), .B(n4720), .C(n2777), .Y(n1996) );
  OAI21X1 U1391 ( .A(n4673), .B(n4720), .C(n2621), .Y(n1997) );
  OAI21X1 U1393 ( .A(n4672), .B(n4720), .C(n2937), .Y(n1998) );
  OAI21X1 U1395 ( .A(n4671), .B(n4720), .C(n2991), .Y(n1999) );
  OAI21X1 U1397 ( .A(n4670), .B(n4720), .C(n2829), .Y(n2000) );
  OAI21X1 U1399 ( .A(n4669), .B(n4720), .C(n2883), .Y(n2001) );
  OAI21X1 U1401 ( .A(n4668), .B(n4720), .C(n2490), .Y(n2002) );
  OAI21X1 U1403 ( .A(n4667), .B(n4720), .C(n2489), .Y(n2003) );
  OAI21X1 U1405 ( .A(n4666), .B(n4720), .C(n2673), .Y(n2004) );
  OAI21X1 U1407 ( .A(n4665), .B(n4720), .C(n2488), .Y(n2005) );
  OAI21X1 U1409 ( .A(n4659), .B(n4720), .C(n2487), .Y(n2006) );
  OAI21X1 U1411 ( .A(n4658), .B(n4720), .C(n2486), .Y(n2007) );
  OAI21X1 U1413 ( .A(n4657), .B(n4720), .C(n2485), .Y(n2008) );
  OAI21X1 U1416 ( .A(n4664), .B(n4718), .C(n3104), .Y(n2009) );
  OAI21X1 U1418 ( .A(n4663), .B(n4719), .C(n3046), .Y(n2010) );
  OAI21X1 U1420 ( .A(n4662), .B(n4718), .C(n3219), .Y(n2011) );
  OAI21X1 U1422 ( .A(n4661), .B(n4719), .C(n3161), .Y(n2012) );
  OAI21X1 U1424 ( .A(n4660), .B(n4718), .C(n3350), .Y(n2013) );
  OAI21X1 U1426 ( .A(n4690), .B(n4719), .C(n3284), .Y(n2014) );
  OAI21X1 U1428 ( .A(n4689), .B(n4718), .C(n3482), .Y(n2015) );
  OAI21X1 U1430 ( .A(n4688), .B(n4719), .C(n3415), .Y(n2016) );
  OAI21X1 U1432 ( .A(n4687), .B(n4718), .C(n2672), .Y(n2017) );
  OAI21X1 U1434 ( .A(n4686), .B(n4719), .C(n3103), .Y(n2018) );
  OAI21X1 U1436 ( .A(n4685), .B(n4718), .C(n2620), .Y(n2019) );
  OAI21X1 U1438 ( .A(n4684), .B(n4719), .C(n2776), .Y(n2020) );
  OAI21X1 U1440 ( .A(n4683), .B(n4718), .C(n2724), .Y(n2021) );
  OAI21X1 U1442 ( .A(n4682), .B(n4718), .C(n3045), .Y(n2022) );
  OAI21X1 U1444 ( .A(n4681), .B(n4719), .C(n3218), .Y(n2023) );
  OAI21X1 U1446 ( .A(n4680), .B(n4719), .C(n3160), .Y(n2024) );
  OAI21X1 U1448 ( .A(n4679), .B(n4718), .C(n3349), .Y(n2025) );
  OAI21X1 U1450 ( .A(n4678), .B(n4719), .C(n3283), .Y(n2026) );
  OAI21X1 U1452 ( .A(n4677), .B(n4718), .C(n3481), .Y(n2027) );
  OAI21X1 U1454 ( .A(n4676), .B(n4719), .C(n3414), .Y(n2028) );
  OAI21X1 U1456 ( .A(n4675), .B(n4718), .C(n2671), .Y(n2029) );
  OAI21X1 U1458 ( .A(n4674), .B(n4718), .C(n2619), .Y(n2030) );
  OAI21X1 U1460 ( .A(n4673), .B(n4718), .C(n2775), .Y(n2031) );
  OAI21X1 U1462 ( .A(n4672), .B(n4718), .C(n2882), .Y(n2032) );
  OAI21X1 U1464 ( .A(n4671), .B(n4718), .C(n2828), .Y(n2033) );
  OAI21X1 U1466 ( .A(n4670), .B(n4718), .C(n2990), .Y(n2034) );
  OAI21X1 U1468 ( .A(n4669), .B(n4718), .C(n2936), .Y(n2035) );
  OAI21X1 U1470 ( .A(n4668), .B(n4718), .C(n2484), .Y(n2036) );
  OAI21X1 U1472 ( .A(n4667), .B(n4718), .C(n2483), .Y(n2037) );
  OAI21X1 U1474 ( .A(n4666), .B(n4718), .C(n2723), .Y(n2038) );
  OAI21X1 U1476 ( .A(n4665), .B(n4718), .C(n2482), .Y(n2039) );
  OAI21X1 U1478 ( .A(n4659), .B(n4718), .C(n2481), .Y(n2040) );
  OAI21X1 U1480 ( .A(n4658), .B(n4718), .C(n2480), .Y(n2041) );
  OAI21X1 U1482 ( .A(n4657), .B(n4718), .C(n2479), .Y(n2042) );
  OAI21X1 U1485 ( .A(n4664), .B(n4716), .C(n3044), .Y(n2043) );
  OAI21X1 U1487 ( .A(n4663), .B(n4717), .C(n3102), .Y(n2044) );
  OAI21X1 U1489 ( .A(n4662), .B(n4716), .C(n3159), .Y(n2045) );
  OAI21X1 U1491 ( .A(n4661), .B(n4717), .C(n3217), .Y(n2046) );
  OAI21X1 U1493 ( .A(n4660), .B(n4716), .C(n3282), .Y(n2047) );
  OAI21X1 U1495 ( .A(n4690), .B(n4717), .C(n3348), .Y(n2048) );
  OAI21X1 U1497 ( .A(n4689), .B(n4716), .C(n3413), .Y(n2049) );
  OAI21X1 U1499 ( .A(n4688), .B(n4717), .C(n3480), .Y(n2050) );
  OAI21X1 U1501 ( .A(n4687), .B(n4716), .C(n2618), .Y(n2051) );
  OAI21X1 U1503 ( .A(n4686), .B(n4717), .C(n3043), .Y(n2052) );
  OAI21X1 U1505 ( .A(n4685), .B(n4716), .C(n2670), .Y(n2053) );
  OAI21X1 U1507 ( .A(n4684), .B(n4717), .C(n2722), .Y(n2054) );
  OAI21X1 U1509 ( .A(n4683), .B(n4716), .C(n2774), .Y(n2055) );
  OAI21X1 U1511 ( .A(n4682), .B(n4716), .C(n3101), .Y(n2056) );
  OAI21X1 U1513 ( .A(n4681), .B(n4717), .C(n3158), .Y(n2057) );
  OAI21X1 U1515 ( .A(n4680), .B(n4717), .C(n3216), .Y(n2058) );
  OAI21X1 U1517 ( .A(n4679), .B(n4716), .C(n3281), .Y(n2059) );
  OAI21X1 U1519 ( .A(n4678), .B(n4717), .C(n3347), .Y(n2060) );
  OAI21X1 U1521 ( .A(n4677), .B(n4716), .C(n3412), .Y(n2061) );
  OAI21X1 U1523 ( .A(n4676), .B(n4717), .C(n3479), .Y(n2062) );
  OAI21X1 U1525 ( .A(n4675), .B(n4716), .C(n2617), .Y(n2063) );
  OAI21X1 U1527 ( .A(n4674), .B(n4716), .C(n2669), .Y(n2064) );
  OAI21X1 U1529 ( .A(n4673), .B(n4716), .C(n2721), .Y(n2065) );
  OAI21X1 U1531 ( .A(n4672), .B(n4716), .C(n2827), .Y(n2066) );
  OAI21X1 U1533 ( .A(n4671), .B(n4716), .C(n2881), .Y(n2067) );
  OAI21X1 U1535 ( .A(n4670), .B(n4716), .C(n2935), .Y(n2068) );
  OAI21X1 U1537 ( .A(n4669), .B(n4716), .C(n2989), .Y(n2069) );
  OAI21X1 U1539 ( .A(n4668), .B(n4716), .C(n2478), .Y(n2070) );
  OAI21X1 U1541 ( .A(n4667), .B(n4716), .C(n2477), .Y(n2071) );
  OAI21X1 U1543 ( .A(n4666), .B(n4716), .C(n2773), .Y(n2072) );
  OAI21X1 U1545 ( .A(n4665), .B(n4716), .C(n2476), .Y(n2073) );
  OAI21X1 U1547 ( .A(n4659), .B(n4716), .C(n2475), .Y(n2074) );
  OAI21X1 U1549 ( .A(n4658), .B(n4716), .C(n2474), .Y(n2075) );
  OAI21X1 U1551 ( .A(n4657), .B(n4716), .C(n2473), .Y(n2076) );
  OAI21X1 U1554 ( .A(n4664), .B(n4714), .C(n2988), .Y(n2077) );
  OAI21X1 U1556 ( .A(n4663), .B(n4715), .C(n2934), .Y(n2078) );
  OAI21X1 U1558 ( .A(n4662), .B(n4714), .C(n2880), .Y(n2079) );
  OAI21X1 U1560 ( .A(n4661), .B(n4715), .C(n2826), .Y(n2080) );
  OAI21X1 U1562 ( .A(n4660), .B(n4714), .C(n2772), .Y(n2081) );
  OAI21X1 U1564 ( .A(n4690), .B(n4715), .C(n2720), .Y(n2082) );
  OAI21X1 U1566 ( .A(n4689), .B(n4714), .C(n2668), .Y(n2083) );
  OAI21X1 U1568 ( .A(n4688), .B(n4715), .C(n2616), .Y(n2084) );
  OAI21X1 U1570 ( .A(n4687), .B(n4714), .C(n3478), .Y(n2085) );
  OAI21X1 U1572 ( .A(n4686), .B(n4715), .C(n2987), .Y(n2086) );
  OAI21X1 U1574 ( .A(n4685), .B(n4714), .C(n3411), .Y(n2087) );
  OAI21X1 U1576 ( .A(n4684), .B(n4715), .C(n3346), .Y(n2088) );
  OAI21X1 U1578 ( .A(n4683), .B(n4714), .C(n3280), .Y(n2089) );
  OAI21X1 U1580 ( .A(n4682), .B(n4714), .C(n2933), .Y(n2090) );
  OAI21X1 U1582 ( .A(n4681), .B(n4715), .C(n2879), .Y(n2091) );
  OAI21X1 U1584 ( .A(n4680), .B(n4715), .C(n2825), .Y(n2092) );
  OAI21X1 U1586 ( .A(n4679), .B(n4714), .C(n2771), .Y(n2093) );
  OAI21X1 U1588 ( .A(n4678), .B(n4715), .C(n2719), .Y(n2094) );
  OAI21X1 U1590 ( .A(n4677), .B(n4714), .C(n2667), .Y(n2095) );
  OAI21X1 U1592 ( .A(n4676), .B(n4715), .C(n2615), .Y(n2096) );
  OAI21X1 U1594 ( .A(n4675), .B(n4714), .C(n3477), .Y(n2097) );
  OAI21X1 U1596 ( .A(n4674), .B(n4714), .C(n3410), .Y(n2098) );
  OAI21X1 U1598 ( .A(n4673), .B(n4714), .C(n3345), .Y(n2099) );
  OAI21X1 U1600 ( .A(n4672), .B(n4714), .C(n3215), .Y(n2100) );
  OAI21X1 U1602 ( .A(n4671), .B(n4714), .C(n3157), .Y(n2101) );
  OAI21X1 U1604 ( .A(n4670), .B(n4714), .C(n3100), .Y(n2102) );
  OAI21X1 U1606 ( .A(n4669), .B(n4714), .C(n3042), .Y(n2103) );
  OAI21X1 U1608 ( .A(n4668), .B(n4714), .C(n2472), .Y(n2104) );
  OAI21X1 U1610 ( .A(n4667), .B(n4714), .C(n2471), .Y(n2105) );
  OAI21X1 U1612 ( .A(n4666), .B(n4714), .C(n3279), .Y(n2106) );
  OAI21X1 U1614 ( .A(n4665), .B(n4714), .C(n2470), .Y(n2107) );
  OAI21X1 U1616 ( .A(n4659), .B(n4714), .C(n2469), .Y(n2108) );
  OAI21X1 U1618 ( .A(n4658), .B(n4714), .C(n2468), .Y(n2109) );
  OAI21X1 U1620 ( .A(n4657), .B(n4714), .C(n2467), .Y(n2110) );
  OAI21X1 U1623 ( .A(n4664), .B(n4712), .C(n2932), .Y(n2111) );
  OAI21X1 U1625 ( .A(n4663), .B(n4713), .C(n2986), .Y(n2112) );
  OAI21X1 U1627 ( .A(n4662), .B(n4712), .C(n2824), .Y(n2113) );
  OAI21X1 U1629 ( .A(n4661), .B(n4713), .C(n2878), .Y(n2114) );
  OAI21X1 U1631 ( .A(n4660), .B(n4712), .C(n2718), .Y(n2115) );
  OAI21X1 U1633 ( .A(n4690), .B(n4713), .C(n2770), .Y(n2116) );
  OAI21X1 U1635 ( .A(n4689), .B(n4712), .C(n2614), .Y(n2117) );
  OAI21X1 U1637 ( .A(n4688), .B(n4713), .C(n2666), .Y(n2118) );
  OAI21X1 U1639 ( .A(n4687), .B(n4712), .C(n3409), .Y(n2119) );
  OAI21X1 U1641 ( .A(n4686), .B(n4713), .C(n2931), .Y(n2120) );
  OAI21X1 U1643 ( .A(n4685), .B(n4712), .C(n3476), .Y(n2121) );
  OAI21X1 U1645 ( .A(n4684), .B(n4713), .C(n3278), .Y(n2122) );
  OAI21X1 U1647 ( .A(n4683), .B(n4712), .C(n3344), .Y(n2123) );
  OAI21X1 U1649 ( .A(n4682), .B(n4712), .C(n2985), .Y(n2124) );
  OAI21X1 U1651 ( .A(n4681), .B(n4713), .C(n2823), .Y(n2125) );
  OAI21X1 U1653 ( .A(n4680), .B(n4713), .C(n2877), .Y(n2126) );
  OAI21X1 U1655 ( .A(n4679), .B(n4712), .C(n2717), .Y(n2127) );
  OAI21X1 U1657 ( .A(n4678), .B(n4713), .C(n2769), .Y(n2128) );
  OAI21X1 U1659 ( .A(n4677), .B(n4712), .C(n2613), .Y(n2129) );
  OAI21X1 U1661 ( .A(n4676), .B(n4713), .C(n2665), .Y(n2130) );
  OAI21X1 U1663 ( .A(n4675), .B(n4712), .C(n3408), .Y(n2131) );
  OAI21X1 U1665 ( .A(n4674), .B(n4712), .C(n3475), .Y(n2132) );
  OAI21X1 U1667 ( .A(n4673), .B(n4712), .C(n3277), .Y(n2133) );
  OAI21X1 U1669 ( .A(n4672), .B(n4712), .C(n3156), .Y(n2134) );
  OAI21X1 U1671 ( .A(n4671), .B(n4712), .C(n3214), .Y(n2135) );
  OAI21X1 U1673 ( .A(n4670), .B(n4712), .C(n3041), .Y(n2136) );
  OAI21X1 U1675 ( .A(n4669), .B(n4712), .C(n3099), .Y(n2137) );
  OAI21X1 U1677 ( .A(n4668), .B(n4712), .C(n2466), .Y(n2138) );
  OAI21X1 U1679 ( .A(n4667), .B(n4712), .C(n2465), .Y(n2139) );
  OAI21X1 U1681 ( .A(n4666), .B(n4712), .C(n3343), .Y(n2140) );
  OAI21X1 U1683 ( .A(n4665), .B(n4712), .C(n2464), .Y(n2141) );
  OAI21X1 U1685 ( .A(n4659), .B(n4712), .C(n1304), .Y(n2142) );
  OAI21X1 U1687 ( .A(n4658), .B(n4712), .C(n153), .Y(n2143) );
  OAI21X1 U1689 ( .A(n4657), .B(n4712), .C(n152), .Y(n2144) );
  OAI21X1 U1692 ( .A(n4664), .B(n4710), .C(n2876), .Y(n2145) );
  OAI21X1 U1694 ( .A(n4663), .B(n4711), .C(n2822), .Y(n2146) );
  OAI21X1 U1696 ( .A(n4662), .B(n4710), .C(n2984), .Y(n2147) );
  OAI21X1 U1698 ( .A(n4661), .B(n4711), .C(n2930), .Y(n2148) );
  OAI21X1 U1700 ( .A(n4660), .B(n4710), .C(n2664), .Y(n2149) );
  OAI21X1 U1702 ( .A(n4690), .B(n4711), .C(n2612), .Y(n2150) );
  OAI21X1 U1704 ( .A(n4689), .B(n4710), .C(n2768), .Y(n2151) );
  OAI21X1 U1706 ( .A(n4688), .B(n4711), .C(n2716), .Y(n2152) );
  OAI21X1 U1708 ( .A(n4687), .B(n4710), .C(n3342), .Y(n2153) );
  OAI21X1 U1710 ( .A(n4686), .B(n4711), .C(n2875), .Y(n2154) );
  OAI21X1 U1712 ( .A(n4685), .B(n4710), .C(n3276), .Y(n2155) );
  OAI21X1 U1714 ( .A(n4684), .B(n4711), .C(n3474), .Y(n2156) );
  OAI21X1 U1716 ( .A(n4683), .B(n4710), .C(n3407), .Y(n2157) );
  OAI21X1 U1718 ( .A(n4682), .B(n4710), .C(n2821), .Y(n2158) );
  OAI21X1 U1720 ( .A(n4681), .B(n4711), .C(n2983), .Y(n2159) );
  OAI21X1 U1722 ( .A(n4680), .B(n4711), .C(n2929), .Y(n2160) );
  OAI21X1 U1724 ( .A(n4679), .B(n4710), .C(n2663), .Y(n2161) );
  OAI21X1 U1726 ( .A(n4678), .B(n4711), .C(n2611), .Y(n2162) );
  OAI21X1 U1728 ( .A(n4677), .B(n4710), .C(n2767), .Y(n2163) );
  OAI21X1 U1730 ( .A(n4676), .B(n4711), .C(n2715), .Y(n2164) );
  OAI21X1 U1732 ( .A(n4675), .B(n4710), .C(n3341), .Y(n2165) );
  OAI21X1 U1734 ( .A(n4674), .B(n4710), .C(n3275), .Y(n2166) );
  OAI21X1 U1736 ( .A(n4673), .B(n4710), .C(n3473), .Y(n2167) );
  OAI21X1 U1738 ( .A(n4672), .B(n4710), .C(n3098), .Y(n2168) );
  OAI21X1 U1740 ( .A(n4671), .B(n4710), .C(n3040), .Y(n2169) );
  OAI21X1 U1742 ( .A(n4670), .B(n4710), .C(n3213), .Y(n2170) );
  OAI21X1 U1744 ( .A(n4669), .B(n4710), .C(n3155), .Y(n2171) );
  OAI21X1 U1746 ( .A(n4668), .B(n4710), .C(n151), .Y(n2172) );
  OAI21X1 U1748 ( .A(n4667), .B(n4710), .C(n150), .Y(n2173) );
  OAI21X1 U1750 ( .A(n4666), .B(n4710), .C(n3406), .Y(n2174) );
  OAI21X1 U1752 ( .A(n4665), .B(n4710), .C(n149), .Y(n2175) );
  OAI21X1 U1754 ( .A(n4659), .B(n4710), .C(n148), .Y(n2176) );
  OAI21X1 U1756 ( .A(n4658), .B(n4710), .C(n147), .Y(n2177) );
  OAI21X1 U1758 ( .A(n4657), .B(n4710), .C(n146), .Y(n2178) );
  NOR3X1 U1761 ( .A(n1288), .B(wr_ptr[3]), .C(n4812), .Y(n759) );
  OAI21X1 U1762 ( .A(n4664), .B(n4708), .C(n2820), .Y(n2179) );
  OAI21X1 U1764 ( .A(n4663), .B(n4708), .C(n2874), .Y(n2180) );
  OAI21X1 U1766 ( .A(n4662), .B(n4709), .C(n2928), .Y(n2181) );
  OAI21X1 U1768 ( .A(n4661), .B(n4708), .C(n2982), .Y(n2182) );
  OAI21X1 U1770 ( .A(n4660), .B(n4709), .C(n2610), .Y(n2183) );
  OAI21X1 U1772 ( .A(n4690), .B(n4708), .C(n2662), .Y(n2184) );
  OAI21X1 U1774 ( .A(n4689), .B(n4709), .C(n2714), .Y(n2185) );
  OAI21X1 U1776 ( .A(n4688), .B(n4708), .C(n2766), .Y(n2186) );
  OAI21X1 U1778 ( .A(n4687), .B(n4709), .C(n3274), .Y(n2187) );
  OAI21X1 U1780 ( .A(n4686), .B(n4708), .C(n2819), .Y(n2188) );
  OAI21X1 U1782 ( .A(n4685), .B(n4709), .C(n3340), .Y(n2189) );
  OAI21X1 U1784 ( .A(n4684), .B(n4708), .C(n3405), .Y(n2190) );
  OAI21X1 U1786 ( .A(n4683), .B(n4709), .C(n3472), .Y(n2191) );
  OAI21X1 U1788 ( .A(n4682), .B(n4709), .C(n2873), .Y(n2192) );
  OAI21X1 U1790 ( .A(n4681), .B(n4708), .C(n2927), .Y(n2193) );
  OAI21X1 U1792 ( .A(n4680), .B(n4708), .C(n2981), .Y(n2194) );
  OAI21X1 U1794 ( .A(n4679), .B(n4709), .C(n2609), .Y(n2195) );
  OAI21X1 U1796 ( .A(n4678), .B(n4708), .C(n2661), .Y(n2196) );
  OAI21X1 U1798 ( .A(n4677), .B(n4709), .C(n2713), .Y(n2197) );
  OAI21X1 U1800 ( .A(n4676), .B(n4708), .C(n2765), .Y(n2198) );
  OAI21X1 U1802 ( .A(n4675), .B(n4708), .C(n3273), .Y(n2199) );
  OAI21X1 U1804 ( .A(n4674), .B(n4708), .C(n3339), .Y(n2200) );
  OAI21X1 U1806 ( .A(n4673), .B(n4709), .C(n3404), .Y(n2201) );
  OAI21X1 U1808 ( .A(n4672), .B(n4708), .C(n3039), .Y(n2202) );
  OAI21X1 U1810 ( .A(n4671), .B(n4708), .C(n3097), .Y(n2203) );
  OAI21X1 U1812 ( .A(n4670), .B(n4708), .C(n3154), .Y(n2204) );
  OAI21X1 U1814 ( .A(n4669), .B(n4708), .C(n3212), .Y(n2205) );
  OAI21X1 U1816 ( .A(n4668), .B(n4708), .C(n145), .Y(n2206) );
  OAI21X1 U1818 ( .A(n4667), .B(n4708), .C(n144), .Y(n2207) );
  OAI21X1 U1820 ( .A(n4666), .B(n4708), .C(n3471), .Y(n2208) );
  OAI21X1 U1822 ( .A(n4665), .B(n4708), .C(n143), .Y(n2209) );
  OAI21X1 U1824 ( .A(n4659), .B(n4708), .C(n142), .Y(n2210) );
  OAI21X1 U1826 ( .A(n4658), .B(n4708), .C(n141), .Y(n2211) );
  OAI21X1 U1828 ( .A(n4657), .B(n4708), .C(n140), .Y(n2212) );
  NOR3X1 U1831 ( .A(wr_ptr[1]), .B(wr_ptr[2]), .C(wr_ptr[0]), .Y(n189) );
  OAI21X1 U1832 ( .A(n4664), .B(n4706), .C(n2764), .Y(n2213) );
  OAI21X1 U1834 ( .A(n4663), .B(n4706), .C(n2712), .Y(n2214) );
  OAI21X1 U1836 ( .A(n4662), .B(n4707), .C(n2660), .Y(n2215) );
  OAI21X1 U1838 ( .A(n4661), .B(n4706), .C(n2608), .Y(n2216) );
  OAI21X1 U1840 ( .A(n4660), .B(n4707), .C(n2980), .Y(n2217) );
  OAI21X1 U1842 ( .A(n4690), .B(n4706), .C(n2926), .Y(n2218) );
  OAI21X1 U1844 ( .A(n4689), .B(n4707), .C(n2872), .Y(n2219) );
  OAI21X1 U1846 ( .A(n4688), .B(n4706), .C(n2818), .Y(n2220) );
  OAI21X1 U1848 ( .A(n4687), .B(n4707), .C(n3211), .Y(n2221) );
  OAI21X1 U1850 ( .A(n4686), .B(n4706), .C(n2763), .Y(n2222) );
  OAI21X1 U1852 ( .A(n4685), .B(n4707), .C(n3153), .Y(n2223) );
  OAI21X1 U1854 ( .A(n4684), .B(n4706), .C(n3096), .Y(n2224) );
  OAI21X1 U1856 ( .A(n4683), .B(n4707), .C(n3038), .Y(n2225) );
  OAI21X1 U1858 ( .A(n4682), .B(n4707), .C(n2711), .Y(n2226) );
  OAI21X1 U1860 ( .A(n4681), .B(n4706), .C(n2659), .Y(n2227) );
  OAI21X1 U1862 ( .A(n4680), .B(n4706), .C(n2607), .Y(n2228) );
  OAI21X1 U1864 ( .A(n4679), .B(n4707), .C(n2979), .Y(n2229) );
  OAI21X1 U1866 ( .A(n4678), .B(n4706), .C(n2925), .Y(n2230) );
  OAI21X1 U1868 ( .A(n4677), .B(n4707), .C(n2871), .Y(n2231) );
  OAI21X1 U1870 ( .A(n4676), .B(n4706), .C(n2817), .Y(n2232) );
  OAI21X1 U1872 ( .A(n4675), .B(n4706), .C(n3210), .Y(n2233) );
  OAI21X1 U1874 ( .A(n4674), .B(n4706), .C(n3152), .Y(n2234) );
  OAI21X1 U1876 ( .A(n4673), .B(n4707), .C(n3095), .Y(n2235) );
  OAI21X1 U1878 ( .A(n4672), .B(n4706), .C(n3470), .Y(n2236) );
  OAI21X1 U1880 ( .A(n4671), .B(n4706), .C(n3403), .Y(n2237) );
  OAI21X1 U1882 ( .A(n4670), .B(n4706), .C(n3338), .Y(n2238) );
  OAI21X1 U1884 ( .A(n4669), .B(n4706), .C(n3272), .Y(n2239) );
  OAI21X1 U1886 ( .A(n4668), .B(n4706), .C(n139), .Y(n2240) );
  OAI21X1 U1888 ( .A(n4667), .B(n4706), .C(n138), .Y(n2241) );
  OAI21X1 U1890 ( .A(n4666), .B(n4706), .C(n3037), .Y(n2242) );
  OAI21X1 U1892 ( .A(n4665), .B(n4706), .C(n137), .Y(n2243) );
  OAI21X1 U1894 ( .A(n4659), .B(n4706), .C(n136), .Y(n2244) );
  OAI21X1 U1896 ( .A(n4658), .B(n4706), .C(n135), .Y(n2245) );
  OAI21X1 U1898 ( .A(n4657), .B(n4706), .C(n134), .Y(n2246) );
  NOR3X1 U1901 ( .A(wr_ptr[1]), .B(wr_ptr[2]), .C(n4808), .Y(n226) );
  OAI21X1 U1902 ( .A(n4664), .B(n4704), .C(n3469), .Y(n2247) );
  OAI21X1 U1904 ( .A(n4663), .B(n4704), .C(n3402), .Y(n2248) );
  OAI21X1 U1906 ( .A(n4662), .B(n4705), .C(n3337), .Y(n2249) );
  OAI21X1 U1908 ( .A(n4661), .B(n4704), .C(n3271), .Y(n2250) );
  OAI21X1 U1910 ( .A(n4660), .B(n4705), .C(n3209), .Y(n2251) );
  OAI21X1 U1912 ( .A(n4690), .B(n4704), .C(n3151), .Y(n2252) );
  OAI21X1 U1914 ( .A(n4689), .B(n4705), .C(n3094), .Y(n2253) );
  OAI21X1 U1916 ( .A(n4688), .B(n4704), .C(n3036), .Y(n2254) );
  OAI21X1 U1918 ( .A(n4687), .B(n4705), .C(n2978), .Y(n2255) );
  OAI21X1 U1920 ( .A(n4686), .B(n4704), .C(n3468), .Y(n2256) );
  OAI21X1 U1922 ( .A(n4685), .B(n4705), .C(n2924), .Y(n2257) );
  OAI21X1 U1924 ( .A(n4684), .B(n4704), .C(n2870), .Y(n2258) );
  OAI21X1 U1926 ( .A(n4683), .B(n4705), .C(n2816), .Y(n2259) );
  OAI21X1 U1928 ( .A(n4682), .B(n4705), .C(n3401), .Y(n2260) );
  OAI21X1 U1930 ( .A(n4681), .B(n4704), .C(n3336), .Y(n2261) );
  OAI21X1 U1932 ( .A(n4680), .B(n4704), .C(n3270), .Y(n2262) );
  OAI21X1 U1934 ( .A(n4679), .B(n4705), .C(n3208), .Y(n2263) );
  OAI21X1 U1936 ( .A(n4678), .B(n4704), .C(n3150), .Y(n2264) );
  OAI21X1 U1938 ( .A(n4677), .B(n4705), .C(n3093), .Y(n2265) );
  OAI21X1 U1940 ( .A(n4676), .B(n4704), .C(n3035), .Y(n2266) );
  OAI21X1 U1942 ( .A(n4675), .B(n4704), .C(n2977), .Y(n2267) );
  OAI21X1 U1944 ( .A(n4674), .B(n4704), .C(n2923), .Y(n2268) );
  OAI21X1 U1946 ( .A(n4673), .B(n4705), .C(n2869), .Y(n2269) );
  OAI21X1 U1948 ( .A(n4672), .B(n4704), .C(n2762), .Y(n2270) );
  OAI21X1 U1950 ( .A(n4671), .B(n4704), .C(n2710), .Y(n2271) );
  OAI21X1 U1952 ( .A(n4670), .B(n4704), .C(n2658), .Y(n2272) );
  OAI21X1 U1954 ( .A(n4669), .B(n4704), .C(n2606), .Y(n2273) );
  OAI21X1 U1956 ( .A(n4668), .B(n4704), .C(n133), .Y(n2274) );
  OAI21X1 U1958 ( .A(n4667), .B(n4704), .C(n132), .Y(n2275) );
  OAI21X1 U1960 ( .A(n4666), .B(n4704), .C(n2815), .Y(n2276) );
  OAI21X1 U1962 ( .A(n4665), .B(n4704), .C(n131), .Y(n2277) );
  OAI21X1 U1964 ( .A(n4659), .B(n4704), .C(n130), .Y(n2278) );
  OAI21X1 U1966 ( .A(n4658), .B(n4704), .C(n129), .Y(n2279) );
  OAI21X1 U1968 ( .A(n4657), .B(n4704), .C(n128), .Y(n2280) );
  NOR3X1 U1971 ( .A(wr_ptr[0]), .B(wr_ptr[2]), .C(n4809), .Y(n262) );
  OAI21X1 U1972 ( .A(n4664), .B(n4702), .C(n3400), .Y(n2281) );
  OAI21X1 U1974 ( .A(n4663), .B(n4702), .C(n3467), .Y(n2282) );
  OAI21X1 U1976 ( .A(n4662), .B(n4703), .C(n3269), .Y(n2283) );
  OAI21X1 U1978 ( .A(n4661), .B(n4702), .C(n3335), .Y(n2284) );
  OAI21X1 U1980 ( .A(n4660), .B(n4703), .C(n3149), .Y(n2285) );
  OAI21X1 U1982 ( .A(n4690), .B(n4702), .C(n3207), .Y(n2286) );
  OAI21X1 U1984 ( .A(n4689), .B(n4703), .C(n3034), .Y(n2287) );
  OAI21X1 U1986 ( .A(n4688), .B(n4702), .C(n3092), .Y(n2288) );
  OAI21X1 U1988 ( .A(n4687), .B(n4703), .C(n2922), .Y(n2289) );
  OAI21X1 U1990 ( .A(n4686), .B(n4702), .C(n3399), .Y(n2290) );
  OAI21X1 U1992 ( .A(n4685), .B(n4703), .C(n2976), .Y(n2291) );
  OAI21X1 U1994 ( .A(n4684), .B(n4702), .C(n2814), .Y(n2292) );
  OAI21X1 U1996 ( .A(n4683), .B(n4703), .C(n2868), .Y(n2293) );
  OAI21X1 U1998 ( .A(n4682), .B(n4703), .C(n3466), .Y(n2294) );
  OAI21X1 U2000 ( .A(n4681), .B(n4702), .C(n3268), .Y(n2295) );
  OAI21X1 U2002 ( .A(n4680), .B(n4702), .C(n3334), .Y(n2296) );
  OAI21X1 U2004 ( .A(n4679), .B(n4703), .C(n3148), .Y(n2297) );
  OAI21X1 U2006 ( .A(n4678), .B(n4702), .C(n3206), .Y(n2298) );
  OAI21X1 U2008 ( .A(n4677), .B(n4703), .C(n3033), .Y(n2299) );
  OAI21X1 U2010 ( .A(n4676), .B(n4702), .C(n3091), .Y(n2300) );
  OAI21X1 U2012 ( .A(n4675), .B(n4702), .C(n2921), .Y(n2301) );
  OAI21X1 U2014 ( .A(n4674), .B(n4702), .C(n2975), .Y(n2302) );
  OAI21X1 U2016 ( .A(n4673), .B(n4703), .C(n2813), .Y(n2303) );
  OAI21X1 U2018 ( .A(n4672), .B(n4702), .C(n2709), .Y(n2304) );
  OAI21X1 U2020 ( .A(n4671), .B(n4702), .C(n2761), .Y(n2305) );
  OAI21X1 U2022 ( .A(n4670), .B(n4702), .C(n2605), .Y(n2306) );
  OAI21X1 U2024 ( .A(n4669), .B(n4702), .C(n2657), .Y(n2307) );
  OAI21X1 U2026 ( .A(n4668), .B(n4702), .C(n127), .Y(n2308) );
  OAI21X1 U2028 ( .A(n4667), .B(n4702), .C(n126), .Y(n2309) );
  OAI21X1 U2030 ( .A(n4666), .B(n4702), .C(n2867), .Y(n2310) );
  OAI21X1 U2032 ( .A(n4665), .B(n4702), .C(n125), .Y(n2311) );
  OAI21X1 U2034 ( .A(n4659), .B(n4702), .C(n124), .Y(n2312) );
  OAI21X1 U2036 ( .A(n4658), .B(n4702), .C(n123), .Y(n2313) );
  OAI21X1 U2038 ( .A(n4657), .B(n4702), .C(n122), .Y(n2314) );
  NOR3X1 U2041 ( .A(n4808), .B(wr_ptr[2]), .C(n4809), .Y(n298) );
  OAI21X1 U2042 ( .A(n4664), .B(n4700), .C(n3333), .Y(n2315) );
  OAI21X1 U2044 ( .A(n4663), .B(n4700), .C(n3267), .Y(n2316) );
  OAI21X1 U2046 ( .A(n4662), .B(n4701), .C(n3465), .Y(n2317) );
  OAI21X1 U2048 ( .A(n4661), .B(n4700), .C(n3398), .Y(n2318) );
  OAI21X1 U2050 ( .A(n4660), .B(n4701), .C(n3090), .Y(n2319) );
  OAI21X1 U2052 ( .A(n4690), .B(n4700), .C(n3032), .Y(n2320) );
  OAI21X1 U2054 ( .A(n4689), .B(n4701), .C(n3205), .Y(n2321) );
  OAI21X1 U2056 ( .A(n4688), .B(n4700), .C(n3147), .Y(n2322) );
  OAI21X1 U2058 ( .A(n4687), .B(n4701), .C(n2866), .Y(n2323) );
  OAI21X1 U2060 ( .A(n4686), .B(n4700), .C(n3332), .Y(n2324) );
  OAI21X1 U2062 ( .A(n4685), .B(n4701), .C(n2812), .Y(n2325) );
  OAI21X1 U2064 ( .A(n4684), .B(n4700), .C(n2974), .Y(n2326) );
  OAI21X1 U2066 ( .A(n4683), .B(n4701), .C(n2920), .Y(n2327) );
  OAI21X1 U2068 ( .A(n4682), .B(n4701), .C(n3266), .Y(n2328) );
  OAI21X1 U2070 ( .A(n4681), .B(n4700), .C(n3464), .Y(n2329) );
  OAI21X1 U2072 ( .A(n4680), .B(n4700), .C(n3397), .Y(n2330) );
  OAI21X1 U2074 ( .A(n4679), .B(n4701), .C(n3089), .Y(n2331) );
  OAI21X1 U2076 ( .A(n4678), .B(n4700), .C(n3031), .Y(n2332) );
  OAI21X1 U2078 ( .A(n4677), .B(n4701), .C(n3204), .Y(n2333) );
  OAI21X1 U2080 ( .A(n4676), .B(n4700), .C(n3146), .Y(n2334) );
  OAI21X1 U2082 ( .A(n4675), .B(n4700), .C(n2865), .Y(n2335) );
  OAI21X1 U2084 ( .A(n4674), .B(n4700), .C(n2811), .Y(n2336) );
  OAI21X1 U2086 ( .A(n4673), .B(n4701), .C(n2973), .Y(n2337) );
  OAI21X1 U2088 ( .A(n4672), .B(n4700), .C(n2656), .Y(n2338) );
  OAI21X1 U2090 ( .A(n4671), .B(n4700), .C(n2604), .Y(n2339) );
  OAI21X1 U2092 ( .A(n4670), .B(n4700), .C(n2760), .Y(n2340) );
  OAI21X1 U2094 ( .A(n4669), .B(n4700), .C(n2708), .Y(n2341) );
  OAI21X1 U2096 ( .A(n4668), .B(n4700), .C(n121), .Y(n2342) );
  OAI21X1 U2098 ( .A(n4667), .B(n4700), .C(n120), .Y(n2343) );
  OAI21X1 U2100 ( .A(n4666), .B(n4700), .C(n2919), .Y(n2344) );
  OAI21X1 U2102 ( .A(n4665), .B(n4700), .C(n119), .Y(n2345) );
  OAI21X1 U2104 ( .A(n4659), .B(n4700), .C(n118), .Y(n2346) );
  OAI21X1 U2106 ( .A(n4658), .B(n4700), .C(n117), .Y(n2347) );
  OAI21X1 U2108 ( .A(n4657), .B(n4700), .C(n116), .Y(n2348) );
  NOR3X1 U2111 ( .A(wr_ptr[0]), .B(wr_ptr[1]), .C(n4810), .Y(n334) );
  OAI21X1 U2112 ( .A(n4664), .B(n4698), .C(n3265), .Y(n2349) );
  OAI21X1 U2114 ( .A(n4663), .B(n4698), .C(n3331), .Y(n2350) );
  OAI21X1 U2116 ( .A(n4662), .B(n4699), .C(n3396), .Y(n2351) );
  OAI21X1 U2118 ( .A(n4661), .B(n4698), .C(n3463), .Y(n2352) );
  OAI21X1 U2120 ( .A(n4660), .B(n4699), .C(n3030), .Y(n2353) );
  OAI21X1 U2122 ( .A(n4690), .B(n4698), .C(n3088), .Y(n2354) );
  OAI21X1 U2124 ( .A(n4689), .B(n4699), .C(n3145), .Y(n2355) );
  OAI21X1 U2126 ( .A(n4688), .B(n4698), .C(n3203), .Y(n2356) );
  OAI21X1 U2128 ( .A(n4687), .B(n4699), .C(n2810), .Y(n2357) );
  OAI21X1 U2130 ( .A(n4686), .B(n4698), .C(n3264), .Y(n2358) );
  OAI21X1 U2132 ( .A(n4685), .B(n4699), .C(n2864), .Y(n2359) );
  OAI21X1 U2134 ( .A(n4684), .B(n4698), .C(n2918), .Y(n2360) );
  OAI21X1 U2136 ( .A(n4683), .B(n4699), .C(n2972), .Y(n2361) );
  OAI21X1 U2138 ( .A(n4682), .B(n4699), .C(n3330), .Y(n2362) );
  OAI21X1 U2140 ( .A(n4681), .B(n4698), .C(n3395), .Y(n2363) );
  OAI21X1 U2142 ( .A(n4680), .B(n4698), .C(n3462), .Y(n2364) );
  OAI21X1 U2144 ( .A(n4679), .B(n4699), .C(n3029), .Y(n2365) );
  OAI21X1 U2146 ( .A(n4678), .B(n4698), .C(n3087), .Y(n2366) );
  OAI21X1 U2148 ( .A(n4677), .B(n4699), .C(n3144), .Y(n2367) );
  OAI21X1 U2150 ( .A(n4676), .B(n4698), .C(n3202), .Y(n2368) );
  OAI21X1 U2152 ( .A(n4675), .B(n4698), .C(n2809), .Y(n2369) );
  OAI21X1 U2154 ( .A(n4674), .B(n4698), .C(n2863), .Y(n2370) );
  OAI21X1 U2156 ( .A(n4673), .B(n4699), .C(n2917), .Y(n2371) );
  OAI21X1 U2158 ( .A(n4672), .B(n4698), .C(n2603), .Y(n2372) );
  OAI21X1 U2160 ( .A(n4671), .B(n4698), .C(n2655), .Y(n2373) );
  OAI21X1 U2162 ( .A(n4670), .B(n4698), .C(n2707), .Y(n2374) );
  OAI21X1 U2164 ( .A(n4669), .B(n4698), .C(n2759), .Y(n2375) );
  OAI21X1 U2166 ( .A(n4668), .B(n4698), .C(n115), .Y(n2376) );
  OAI21X1 U2168 ( .A(n4667), .B(n4698), .C(n114), .Y(n2377) );
  OAI21X1 U2170 ( .A(n4666), .B(n4698), .C(n2971), .Y(n2378) );
  OAI21X1 U2172 ( .A(n4665), .B(n4698), .C(n113), .Y(n2379) );
  OAI21X1 U2174 ( .A(n4659), .B(n4698), .C(n112), .Y(n2380) );
  OAI21X1 U2176 ( .A(n4658), .B(n4698), .C(n111), .Y(n2381) );
  OAI21X1 U2178 ( .A(n4657), .B(n4698), .C(n110), .Y(n2382) );
  NOR3X1 U2181 ( .A(n4808), .B(wr_ptr[1]), .C(n4810), .Y(n370) );
  OAI21X1 U2182 ( .A(n4664), .B(n4696), .C(n3201), .Y(n2383) );
  OAI21X1 U2184 ( .A(n4663), .B(n4696), .C(n3143), .Y(n2384) );
  OAI21X1 U2186 ( .A(n4662), .B(n4697), .C(n3086), .Y(n2385) );
  OAI21X1 U2188 ( .A(n4661), .B(n4696), .C(n3028), .Y(n2386) );
  OAI21X1 U2190 ( .A(n4660), .B(n4697), .C(n3461), .Y(n2387) );
  OAI21X1 U2192 ( .A(n4690), .B(n4696), .C(n3394), .Y(n2388) );
  OAI21X1 U2194 ( .A(n4689), .B(n4697), .C(n3329), .Y(n2389) );
  OAI21X1 U2196 ( .A(n4688), .B(n4696), .C(n3263), .Y(n2390) );
  OAI21X1 U2198 ( .A(n4687), .B(n4697), .C(n2758), .Y(n2391) );
  OAI21X1 U2200 ( .A(n4686), .B(n4696), .C(n3200), .Y(n2392) );
  OAI21X1 U2202 ( .A(n4685), .B(n4697), .C(n2706), .Y(n2393) );
  OAI21X1 U2204 ( .A(n4684), .B(n4696), .C(n2654), .Y(n2394) );
  OAI21X1 U2206 ( .A(n4683), .B(n4697), .C(n2602), .Y(n2395) );
  OAI21X1 U2208 ( .A(n4682), .B(n4697), .C(n3142), .Y(n2396) );
  OAI21X1 U2210 ( .A(n4681), .B(n4696), .C(n3085), .Y(n2397) );
  OAI21X1 U2212 ( .A(n4680), .B(n4696), .C(n3027), .Y(n2398) );
  OAI21X1 U2214 ( .A(n4679), .B(n4697), .C(n3460), .Y(n2399) );
  OAI21X1 U2216 ( .A(n4678), .B(n4696), .C(n3393), .Y(n2400) );
  OAI21X1 U2218 ( .A(n4677), .B(n4697), .C(n3328), .Y(n2401) );
  OAI21X1 U2220 ( .A(n4676), .B(n4696), .C(n3262), .Y(n2402) );
  OAI21X1 U2222 ( .A(n4675), .B(n4696), .C(n2757), .Y(n2403) );
  OAI21X1 U2224 ( .A(n4674), .B(n4696), .C(n2705), .Y(n2404) );
  OAI21X1 U2226 ( .A(n4673), .B(n4697), .C(n2653), .Y(n2405) );
  OAI21X1 U2228 ( .A(n4672), .B(n4696), .C(n2970), .Y(n2406) );
  OAI21X1 U2230 ( .A(n4671), .B(n4696), .C(n2916), .Y(n2407) );
  OAI21X1 U2232 ( .A(n4670), .B(n4696), .C(n2862), .Y(n2408) );
  OAI21X1 U2234 ( .A(n4669), .B(n4696), .C(n2808), .Y(n2409) );
  OAI21X1 U2236 ( .A(n4668), .B(n4696), .C(n109), .Y(n2410) );
  OAI21X1 U2238 ( .A(n4667), .B(n4696), .C(n108), .Y(n2411) );
  OAI21X1 U2240 ( .A(n4666), .B(n4696), .C(n2601), .Y(n2412) );
  OAI21X1 U2242 ( .A(n4665), .B(n4696), .C(n107), .Y(n2413) );
  OAI21X1 U2244 ( .A(n4659), .B(n4696), .C(n106), .Y(n2414) );
  OAI21X1 U2246 ( .A(n4658), .B(n4696), .C(n105), .Y(n2415) );
  OAI21X1 U2248 ( .A(n4657), .B(n4696), .C(n104), .Y(n2416) );
  NOR3X1 U2251 ( .A(n4809), .B(wr_ptr[0]), .C(n4810), .Y(n406) );
  OAI21X1 U2252 ( .A(n4664), .B(n4694), .C(n3141), .Y(n2417) );
  OAI21X1 U2254 ( .A(n4663), .B(n4694), .C(n3199), .Y(n2418) );
  OAI21X1 U2256 ( .A(n4662), .B(n4695), .C(n3026), .Y(n2419) );
  OAI21X1 U2258 ( .A(n4661), .B(n4694), .C(n3084), .Y(n2420) );
  OAI21X1 U2260 ( .A(n4660), .B(n4695), .C(n3392), .Y(n2421) );
  OAI21X1 U2262 ( .A(n4690), .B(n4694), .C(n3459), .Y(n2422) );
  OAI21X1 U2264 ( .A(n4689), .B(n4695), .C(n3261), .Y(n2423) );
  OAI21X1 U2266 ( .A(n4688), .B(n4694), .C(n3327), .Y(n2424) );
  OAI21X1 U2268 ( .A(n4687), .B(n4695), .C(n2704), .Y(n2425) );
  OAI21X1 U2270 ( .A(n4686), .B(n4694), .C(n3140), .Y(n2426) );
  OAI21X1 U2272 ( .A(n4685), .B(n4695), .C(n2756), .Y(n2427) );
  OAI21X1 U2274 ( .A(n4684), .B(n4694), .C(n2600), .Y(n2428) );
  OAI21X1 U2276 ( .A(n4683), .B(n4695), .C(n2652), .Y(n2429) );
  OAI21X1 U2278 ( .A(n4682), .B(n4695), .C(n3198), .Y(n2430) );
  OAI21X1 U2280 ( .A(n4681), .B(n4694), .C(n3025), .Y(n2431) );
  OAI21X1 U2282 ( .A(n4680), .B(n4694), .C(n3083), .Y(n2432) );
  OAI21X1 U2284 ( .A(n4679), .B(n4695), .C(n3391), .Y(n2433) );
  OAI21X1 U2286 ( .A(n4678), .B(n4694), .C(n3458), .Y(n2434) );
  OAI21X1 U2288 ( .A(n4677), .B(n4695), .C(n3260), .Y(n2435) );
  OAI21X1 U2290 ( .A(n4676), .B(n4694), .C(n3326), .Y(n2436) );
  OAI21X1 U2292 ( .A(n4675), .B(n4694), .C(n2703), .Y(n2437) );
  OAI21X1 U2294 ( .A(n4674), .B(n4694), .C(n2755), .Y(n2438) );
  OAI21X1 U2296 ( .A(n4673), .B(n4695), .C(n2599), .Y(n2439) );
  OAI21X1 U2298 ( .A(n4672), .B(n4694), .C(n2915), .Y(n2440) );
  OAI21X1 U2300 ( .A(n4671), .B(n4694), .C(n2969), .Y(n2441) );
  OAI21X1 U2302 ( .A(n4670), .B(n4694), .C(n2807), .Y(n2442) );
  OAI21X1 U2304 ( .A(n4669), .B(n4694), .C(n2861), .Y(n2443) );
  OAI21X1 U2306 ( .A(n4668), .B(n4694), .C(n103), .Y(n2444) );
  OAI21X1 U2308 ( .A(n4667), .B(n4694), .C(n102), .Y(n2445) );
  OAI21X1 U2310 ( .A(n4666), .B(n4694), .C(n2651), .Y(n2446) );
  OAI21X1 U2312 ( .A(n4665), .B(n4694), .C(n101), .Y(n2447) );
  OAI21X1 U2314 ( .A(n4659), .B(n4694), .C(n94), .Y(n2448) );
  OAI21X1 U2316 ( .A(n4658), .B(n4694), .C(n93), .Y(n2449) );
  OAI21X1 U2318 ( .A(n4657), .B(n4694), .C(n92), .Y(n2450) );
  NOR3X1 U2321 ( .A(n4809), .B(n4808), .C(n4810), .Y(n442) );
  NOR3X1 U2322 ( .A(n4811), .B(n1288), .C(n4812), .Y(n1040) );
  OAI21X1 U2323 ( .A(n4812), .B(n3524), .C(n3259), .Y(n2451) );
  OAI21X1 U2325 ( .A(n4811), .B(n3524), .C(n3197), .Y(n2452) );
  OAI21X1 U2327 ( .A(n4810), .B(n3524), .C(n3139), .Y(n2453) );
  OAI21X1 U2329 ( .A(n4809), .B(n3524), .C(n3081), .Y(n2454) );
  OAI21X1 U2331 ( .A(n4808), .B(n3524), .C(n3023), .Y(n2455) );
  OAI21X1 U2335 ( .A(n1295), .B(n4813), .C(n3082), .Y(n2456) );
  AOI22X1 U2336 ( .A(n99), .B(n1297), .C(n87), .D(n1298), .Y(n1296) );
  OAI21X1 U2337 ( .A(n1295), .B(n4763), .C(n3254), .Y(n2457) );
  AOI22X1 U2338 ( .A(n98), .B(n1297), .C(n86), .D(n1298), .Y(n1299) );
  OAI21X1 U2339 ( .A(n1295), .B(n4764), .C(n3196), .Y(n2458) );
  AOI22X1 U2340 ( .A(n97), .B(n1297), .C(n85), .D(n1298), .Y(n1300) );
  OAI21X1 U2341 ( .A(n1295), .B(n4814), .C(n3322), .Y(n2459) );
  AOI22X1 U2342 ( .A(n96), .B(n1297), .C(n84), .D(n1298), .Y(n1301) );
  OAI21X1 U2343 ( .A(n1295), .B(n95), .C(n3024), .Y(n2460) );
  AOI22X1 U2344 ( .A(n95), .B(n1297), .C(n95), .D(n1298), .Y(n1302) );
  AOI22X1 U2345 ( .A(n76), .B(n4691), .C(n23), .D(n1305), .Y(n1303) );
  AOI22X1 U2346 ( .A(n75), .B(n4691), .C(n22), .D(n1305), .Y(n1306) );
  AOI22X1 U2347 ( .A(n74), .B(n4693), .C(n21), .D(n1305), .Y(n1307) );
  AOI22X1 U2348 ( .A(n73), .B(n4693), .C(n20), .D(n1305), .Y(n1308) );
  AOI22X1 U2349 ( .A(n4585), .B(n4693), .C(n4592), .D(n1305), .Y(n1309) );
  AOI22X1 U2350 ( .A(data_out[33]), .B(n4692), .C(n24), .D(n4693), .Y(n1310)
         );
  AOI22X1 U2351 ( .A(data_out[32]), .B(n4692), .C(n25), .D(n4691), .Y(n1311)
         );
  AOI22X1 U2352 ( .A(data_out[31]), .B(n4692), .C(n26), .D(n4691), .Y(n1312)
         );
  AOI22X1 U2353 ( .A(data_out[30]), .B(n4692), .C(n27), .D(n4693), .Y(n1313)
         );
  AOI22X1 U2354 ( .A(data_out[29]), .B(n4692), .C(n28), .D(n4691), .Y(n1314)
         );
  AOI22X1 U2355 ( .A(data_out[28]), .B(n4692), .C(n29), .D(n4693), .Y(n1315)
         );
  AOI22X1 U2356 ( .A(data_out[27]), .B(n4692), .C(n30), .D(n4691), .Y(n1316)
         );
  AOI22X1 U2357 ( .A(data_out[26]), .B(n4692), .C(n31), .D(n4691), .Y(n1317)
         );
  AOI22X1 U2358 ( .A(data_out[25]), .B(n4692), .C(n32), .D(n4693), .Y(n1318)
         );
  AOI22X1 U2359 ( .A(data_out[24]), .B(n4692), .C(n33), .D(n4691), .Y(n1319)
         );
  AOI22X1 U2360 ( .A(data_out[23]), .B(n4692), .C(n34), .D(n4691), .Y(n1320)
         );
  AOI22X1 U2361 ( .A(data_out[22]), .B(n4692), .C(n35), .D(n4691), .Y(n1321)
         );
  AOI22X1 U2362 ( .A(data_out[21]), .B(n4692), .C(n36), .D(n4691), .Y(n1322)
         );
  AOI22X1 U2363 ( .A(data_out[20]), .B(n4692), .C(n37), .D(n4691), .Y(n1323)
         );
  AOI22X1 U2364 ( .A(data_out[19]), .B(n4692), .C(n38), .D(n4691), .Y(n1324)
         );
  AOI22X1 U2365 ( .A(data_out[18]), .B(n3525), .C(n39), .D(n4691), .Y(n1325)
         );
  AOI22X1 U2366 ( .A(data_out[17]), .B(n3525), .C(n40), .D(n4691), .Y(n1326)
         );
  AOI22X1 U2367 ( .A(data_out[16]), .B(n3525), .C(n41), .D(n4691), .Y(n1327)
         );
  AOI22X1 U2368 ( .A(data_out[15]), .B(n3525), .C(n42), .D(n4691), .Y(n1328)
         );
  AOI22X1 U2369 ( .A(data_out[14]), .B(n3525), .C(n43), .D(n4691), .Y(n1329)
         );
  AOI22X1 U2370 ( .A(data_out[13]), .B(n3525), .C(n44), .D(n4691), .Y(n1330)
         );
  AOI22X1 U2371 ( .A(data_out[12]), .B(n3525), .C(n45), .D(n4691), .Y(n1331)
         );
  AOI22X1 U2372 ( .A(data_out[11]), .B(n3525), .C(n46), .D(n4691), .Y(n1332)
         );
  AOI22X1 U2373 ( .A(data_out[10]), .B(n3525), .C(n47), .D(n4693), .Y(n1333)
         );
  AOI22X1 U2374 ( .A(data_out[9]), .B(n4692), .C(n48), .D(n4693), .Y(n1334) );
  AOI22X1 U2375 ( .A(data_out[8]), .B(n4692), .C(n49), .D(n4691), .Y(n1335) );
  AOI22X1 U2376 ( .A(data_out[7]), .B(n4692), .C(n50), .D(n4691), .Y(n1336) );
  AOI22X1 U2377 ( .A(data_out[6]), .B(n4692), .C(n51), .D(n4691), .Y(n1337) );
  AOI22X1 U2378 ( .A(data_out[5]), .B(n4692), .C(n52), .D(n4691), .Y(n1338) );
  AOI22X1 U2379 ( .A(data_out[4]), .B(n4692), .C(n53), .D(n4691), .Y(n1339) );
  AOI22X1 U2380 ( .A(data_out[3]), .B(n3525), .C(n54), .D(n4693), .Y(n1340) );
  AOI22X1 U2381 ( .A(data_out[2]), .B(n4692), .C(n55), .D(n4691), .Y(n1341) );
  AOI22X1 U2382 ( .A(data_out[1]), .B(n4692), .C(n56), .D(n4693), .Y(n1342) );
  AOI22X1 U2383 ( .A(data_out[0]), .B(n4692), .C(n57), .D(n4691), .Y(n1343) );
  OAI21X1 U2385 ( .A(n3324), .B(n4807), .C(n3323), .Y(n2461) );
  NAND3X1 U2387 ( .A(n3325), .B(n4758), .C(n3390), .Y(n1346) );
  NAND3X1 U2388 ( .A(n1350), .B(n4765), .C(n1351), .Y(n1349) );
  NOR3X1 U2389 ( .A(n3520), .B(fillcount[3]), .C(fillcount[2]), .Y(n1351) );
  OAI21X1 U2391 ( .A(n1295), .B(n4806), .C(n3388), .Y(n2462) );
  AOI22X1 U2392 ( .A(n100), .B(n1297), .C(n88), .D(n1298), .Y(n1353) );
  OAI21X1 U2394 ( .A(n3257), .B(n4805), .C(n3256), .Y(n2463) );
  NAND3X1 U2396 ( .A(n3258), .B(n4758), .C(n3523), .Y(n1356) );
  NAND3X1 U2397 ( .A(get), .B(n4807), .C(n1355), .Y(n1344) );
  NAND3X1 U2398 ( .A(n3389), .B(n1293), .C(n1361), .Y(n1358) );
  NOR3X1 U2399 ( .A(n3453), .B(fillcount[5]), .C(n4813), .Y(n1361) );
  NAND3X1 U2402 ( .A(n1359), .B(n4807), .C(get), .Y(n1345) );
  HAX1 add_45_U1_1_1 ( .A(fillcount[1]), .B(fillcount[0]), .YC(add_45_carry[2]), .YS(n84) );
  HAX1 add_45_U1_1_2 ( .A(fillcount[2]), .B(add_45_carry[2]), .YC(
        add_45_carry[3]), .YS(n85) );
  HAX1 add_45_U1_1_3 ( .A(fillcount[3]), .B(add_45_carry[3]), .YC(
        add_45_carry[4]), .YS(n86) );
  HAX1 add_45_U1_1_4 ( .A(fillcount[4]), .B(add_45_carry[4]), .YC(
        add_45_carry[5]), .YS(n87) );
  HAX1 r308_U1_1_1 ( .A(n20), .B(n4591), .YC(r308_carry[2]), .YS(n73) );
  HAX1 r308_U1_1_2 ( .A(n21), .B(r308_carry[2]), .YC(r308_carry[3]), .YS(n74)
         );
  HAX1 r308_U1_1_3 ( .A(n22), .B(r308_carry[3]), .YC(r308_carry[4]), .YS(n75)
         );
  HAX1 r307_U1_1_1 ( .A(wr_ptr[1]), .B(wr_ptr[0]), .YC(r307_carry[2]), .YS(n68) );
  HAX1 r307_U1_1_2 ( .A(wr_ptr[2]), .B(r307_carry[2]), .YC(r307_carry[3]), 
        .YS(n69) );
  HAX1 r307_U1_1_3 ( .A(wr_ptr[3]), .B(r307_carry[3]), .YC(r307_carry[4]), 
        .YS(n70) );
  OR2X1 U3 ( .A(n3255), .B(reset), .Y(n1294) );
  OR2X1 U4 ( .A(n3456), .B(n1293), .Y(n1295) );
  OR2X1 U5 ( .A(n3522), .B(fillcount[4]), .Y(n4762) );
  AND2X1 U6 ( .A(n3324), .B(n3456), .Y(n1347) );
  AND2X1 U7 ( .A(n1293), .B(n3257), .Y(n1357) );
  AND2X1 U8 ( .A(n3390), .B(n1294), .Y(n1288) );
  AND2X1 U9 ( .A(n1354), .B(n3255), .Y(n1293) );
  AND2X1 U10 ( .A(n1294), .B(n3523), .Y(n3525) );
  BUFX2 U11 ( .A(n1343), .Y(n1) );
  BUFX2 U12 ( .A(n1342), .Y(n2) );
  BUFX2 U13 ( .A(n1341), .Y(n3) );
  BUFX2 U14 ( .A(n1340), .Y(n4) );
  BUFX2 U15 ( .A(n1339), .Y(n5) );
  BUFX2 U16 ( .A(n1338), .Y(n6) );
  BUFX2 U17 ( .A(n1337), .Y(n7) );
  BUFX2 U18 ( .A(n1336), .Y(n8) );
  BUFX2 U19 ( .A(n1335), .Y(n9) );
  BUFX2 U20 ( .A(n1334), .Y(n10) );
  BUFX2 U21 ( .A(n1333), .Y(n11) );
  BUFX2 U22 ( .A(n1332), .Y(n12) );
  BUFX2 U23 ( .A(n1331), .Y(n13) );
  BUFX2 U24 ( .A(n1330), .Y(n14) );
  BUFX2 U25 ( .A(n1329), .Y(n15) );
  BUFX2 U26 ( .A(n1328), .Y(n16) );
  BUFX2 U27 ( .A(n1327), .Y(n17) );
  BUFX2 U28 ( .A(n1326), .Y(n18) );
  BUFX2 U29 ( .A(n1325), .Y(n58) );
  BUFX2 U30 ( .A(n1324), .Y(n59) );
  BUFX2 U31 ( .A(n1323), .Y(n60) );
  BUFX2 U32 ( .A(n1322), .Y(n61) );
  BUFX2 U33 ( .A(n1321), .Y(n62) );
  BUFX2 U34 ( .A(n1320), .Y(n63) );
  BUFX2 U35 ( .A(n1319), .Y(n64) );
  BUFX2 U36 ( .A(n1318), .Y(n65) );
  BUFX2 U37 ( .A(n1317), .Y(n66) );
  BUFX2 U38 ( .A(n1316), .Y(n67) );
  BUFX2 U39 ( .A(n1315), .Y(n72) );
  BUFX2 U40 ( .A(n1314), .Y(n77) );
  BUFX2 U41 ( .A(n1313), .Y(n78) );
  BUFX2 U42 ( .A(n1312), .Y(n79) );
  BUFX2 U43 ( .A(n1311), .Y(n80) );
  BUFX2 U44 ( .A(n1310), .Y(n81) );
  BUFX2 U45 ( .A(n1309), .Y(n82) );
  BUFX2 U46 ( .A(n1308), .Y(n83) );
  BUFX2 U47 ( .A(n1307), .Y(n89) );
  BUFX2 U48 ( .A(n1306), .Y(n90) );
  BUFX2 U49 ( .A(n1303), .Y(n91) );
  AND2X1 U50 ( .A(n1040), .B(n442), .Y(n1251) );
  AND2X1 U51 ( .A(n1040), .B(n406), .Y(n1216) );
  AND2X1 U52 ( .A(n1040), .B(n370), .Y(n1181) );
  AND2X1 U53 ( .A(n1040), .B(n334), .Y(n1146) );
  AND2X1 U54 ( .A(n1040), .B(n298), .Y(n1111) );
  AND2X1 U55 ( .A(n1040), .B(n262), .Y(n1076) );
  AND2X1 U56 ( .A(n1040), .B(n226), .Y(n1041) );
  AND2X1 U57 ( .A(n1040), .B(n189), .Y(n1005) );
  AND2X1 U58 ( .A(n759), .B(n442), .Y(n970) );
  AND2X1 U59 ( .A(n759), .B(n406), .Y(n935) );
  AND2X1 U60 ( .A(n759), .B(n370), .Y(n900) );
  AND2X1 U61 ( .A(n759), .B(n334), .Y(n865) );
  AND2X1 U62 ( .A(n759), .B(n298), .Y(n830) );
  AND2X1 U63 ( .A(n759), .B(n262), .Y(n795) );
  AND2X1 U64 ( .A(n759), .B(n226), .Y(n760) );
  AND2X1 U65 ( .A(n759), .B(n189), .Y(n724) );
  AND2X1 U66 ( .A(n478), .B(n442), .Y(n689) );
  AND2X1 U67 ( .A(n478), .B(n406), .Y(n654) );
  AND2X1 U68 ( .A(n478), .B(n370), .Y(n619) );
  AND2X1 U69 ( .A(n478), .B(n334), .Y(n584) );
  AND2X1 U70 ( .A(n478), .B(n298), .Y(n549) );
  AND2X1 U71 ( .A(n478), .B(n262), .Y(n514) );
  AND2X1 U72 ( .A(n478), .B(n226), .Y(n479) );
  AND2X1 U73 ( .A(n478), .B(n189), .Y(n443) );
  AND2X1 U74 ( .A(n442), .B(n190), .Y(n407) );
  AND2X1 U75 ( .A(n406), .B(n190), .Y(n371) );
  AND2X1 U76 ( .A(n370), .B(n190), .Y(n335) );
  AND2X1 U77 ( .A(n334), .B(n190), .Y(n299) );
  AND2X1 U78 ( .A(n298), .B(n190), .Y(n263) );
  AND2X1 U79 ( .A(n262), .B(n190), .Y(n227) );
  AND2X1 U80 ( .A(n226), .B(n190), .Y(n191) );
  AND2X1 U81 ( .A(n189), .B(n190), .Y(n154) );
  AND2X1 U82 ( .A(fifo_array[1087]), .B(n4694), .Y(n1285) );
  INVX1 U83 ( .A(n1285), .Y(n92) );
  AND2X1 U84 ( .A(fifo_array[1086]), .B(n4695), .Y(n1284) );
  INVX1 U85 ( .A(n1284), .Y(n93) );
  AND2X1 U86 ( .A(fifo_array[1085]), .B(n4694), .Y(n1283) );
  INVX1 U87 ( .A(n1283), .Y(n94) );
  AND2X1 U88 ( .A(fifo_array[1084]), .B(n4695), .Y(n1282) );
  INVX1 U89 ( .A(n1282), .Y(n101) );
  AND2X1 U90 ( .A(fifo_array[1082]), .B(n4695), .Y(n1280) );
  INVX1 U91 ( .A(n1280), .Y(n102) );
  AND2X1 U92 ( .A(fifo_array[1081]), .B(n4695), .Y(n1279) );
  INVX1 U93 ( .A(n1279), .Y(n103) );
  AND2X1 U94 ( .A(fifo_array[1053]), .B(n4696), .Y(n1250) );
  INVX1 U95 ( .A(n1250), .Y(n104) );
  AND2X1 U96 ( .A(fifo_array[1052]), .B(n4697), .Y(n1249) );
  INVX1 U97 ( .A(n1249), .Y(n105) );
  AND2X1 U98 ( .A(fifo_array[1051]), .B(n4696), .Y(n1248) );
  INVX1 U99 ( .A(n1248), .Y(n106) );
  AND2X1 U100 ( .A(fifo_array[1050]), .B(n4697), .Y(n1247) );
  INVX1 U101 ( .A(n1247), .Y(n107) );
  AND2X1 U102 ( .A(fifo_array[1048]), .B(n4697), .Y(n1245) );
  INVX1 U104 ( .A(n1245), .Y(n108) );
  AND2X1 U106 ( .A(fifo_array[1047]), .B(n4697), .Y(n1244) );
  INVX1 U108 ( .A(n1244), .Y(n109) );
  AND2X1 U110 ( .A(fifo_array[1019]), .B(n4698), .Y(n1215) );
  INVX1 U112 ( .A(n1215), .Y(n110) );
  AND2X1 U114 ( .A(fifo_array[1018]), .B(n4699), .Y(n1214) );
  INVX1 U116 ( .A(n1214), .Y(n111) );
  AND2X1 U118 ( .A(fifo_array[1017]), .B(n4698), .Y(n1213) );
  INVX1 U120 ( .A(n1213), .Y(n112) );
  AND2X1 U122 ( .A(fifo_array[1016]), .B(n4699), .Y(n1212) );
  INVX1 U124 ( .A(n1212), .Y(n113) );
  AND2X1 U126 ( .A(fifo_array[1014]), .B(n4699), .Y(n1210) );
  INVX1 U128 ( .A(n1210), .Y(n114) );
  AND2X1 U130 ( .A(fifo_array[1013]), .B(n4699), .Y(n1209) );
  INVX1 U132 ( .A(n1209), .Y(n115) );
  AND2X1 U134 ( .A(fifo_array[985]), .B(n4700), .Y(n1180) );
  INVX1 U136 ( .A(n1180), .Y(n116) );
  AND2X1 U138 ( .A(fifo_array[984]), .B(n4701), .Y(n1179) );
  INVX1 U140 ( .A(n1179), .Y(n117) );
  AND2X1 U142 ( .A(fifo_array[983]), .B(n4700), .Y(n1178) );
  INVX1 U144 ( .A(n1178), .Y(n118) );
  AND2X1 U146 ( .A(fifo_array[982]), .B(n4701), .Y(n1177) );
  INVX1 U148 ( .A(n1177), .Y(n119) );
  AND2X1 U150 ( .A(fifo_array[980]), .B(n4701), .Y(n1175) );
  INVX1 U152 ( .A(n1175), .Y(n120) );
  AND2X1 U154 ( .A(fifo_array[979]), .B(n4701), .Y(n1174) );
  INVX1 U156 ( .A(n1174), .Y(n121) );
  AND2X1 U158 ( .A(fifo_array[951]), .B(n4702), .Y(n1145) );
  INVX1 U160 ( .A(n1145), .Y(n122) );
  AND2X1 U162 ( .A(fifo_array[950]), .B(n4703), .Y(n1144) );
  INVX1 U164 ( .A(n1144), .Y(n123) );
  AND2X1 U166 ( .A(fifo_array[949]), .B(n4702), .Y(n1143) );
  INVX1 U168 ( .A(n1143), .Y(n124) );
  AND2X1 U170 ( .A(fifo_array[948]), .B(n4703), .Y(n1142) );
  INVX1 U171 ( .A(n1142), .Y(n125) );
  AND2X1 U173 ( .A(fifo_array[946]), .B(n4703), .Y(n1140) );
  INVX1 U175 ( .A(n1140), .Y(n126) );
  AND2X1 U177 ( .A(fifo_array[945]), .B(n4703), .Y(n1139) );
  INVX1 U179 ( .A(n1139), .Y(n127) );
  AND2X1 U181 ( .A(fifo_array[917]), .B(n4704), .Y(n1110) );
  INVX1 U183 ( .A(n1110), .Y(n128) );
  AND2X1 U185 ( .A(fifo_array[916]), .B(n4705), .Y(n1109) );
  INVX1 U187 ( .A(n1109), .Y(n129) );
  AND2X1 U189 ( .A(fifo_array[915]), .B(n4704), .Y(n1108) );
  INVX1 U191 ( .A(n1108), .Y(n130) );
  AND2X1 U193 ( .A(fifo_array[914]), .B(n4705), .Y(n1107) );
  INVX1 U195 ( .A(n1107), .Y(n131) );
  AND2X1 U197 ( .A(fifo_array[912]), .B(n4705), .Y(n1105) );
  INVX1 U199 ( .A(n1105), .Y(n132) );
  AND2X1 U201 ( .A(fifo_array[911]), .B(n4705), .Y(n1104) );
  INVX1 U203 ( .A(n1104), .Y(n133) );
  AND2X1 U205 ( .A(fifo_array[883]), .B(n4706), .Y(n1075) );
  INVX1 U207 ( .A(n1075), .Y(n134) );
  AND2X1 U209 ( .A(fifo_array[882]), .B(n4707), .Y(n1074) );
  INVX1 U211 ( .A(n1074), .Y(n135) );
  AND2X1 U213 ( .A(fifo_array[881]), .B(n4706), .Y(n1073) );
  INVX1 U215 ( .A(n1073), .Y(n136) );
  AND2X1 U217 ( .A(fifo_array[880]), .B(n4707), .Y(n1072) );
  INVX1 U219 ( .A(n1072), .Y(n137) );
  AND2X1 U221 ( .A(fifo_array[878]), .B(n4707), .Y(n1070) );
  INVX1 U223 ( .A(n1070), .Y(n138) );
  AND2X1 U225 ( .A(fifo_array[877]), .B(n4707), .Y(n1069) );
  INVX1 U227 ( .A(n1069), .Y(n139) );
  AND2X1 U229 ( .A(fifo_array[849]), .B(n4708), .Y(n1039) );
  INVX1 U231 ( .A(n1039), .Y(n140) );
  AND2X1 U233 ( .A(fifo_array[848]), .B(n4709), .Y(n1038) );
  INVX1 U235 ( .A(n1038), .Y(n141) );
  AND2X1 U237 ( .A(fifo_array[847]), .B(n4708), .Y(n1037) );
  INVX1 U239 ( .A(n1037), .Y(n142) );
  AND2X1 U240 ( .A(fifo_array[846]), .B(n4709), .Y(n1036) );
  INVX1 U242 ( .A(n1036), .Y(n143) );
  AND2X1 U244 ( .A(fifo_array[844]), .B(n4709), .Y(n1034) );
  INVX1 U246 ( .A(n1034), .Y(n144) );
  AND2X1 U248 ( .A(fifo_array[843]), .B(n4709), .Y(n1033) );
  INVX1 U250 ( .A(n1033), .Y(n145) );
  AND2X1 U252 ( .A(fifo_array[815]), .B(n4711), .Y(n1004) );
  INVX1 U254 ( .A(n1004), .Y(n146) );
  AND2X1 U256 ( .A(fifo_array[814]), .B(n4711), .Y(n1003) );
  INVX1 U258 ( .A(n1003), .Y(n147) );
  AND2X1 U260 ( .A(fifo_array[813]), .B(n4711), .Y(n1002) );
  INVX1 U262 ( .A(n1002), .Y(n148) );
  AND2X1 U264 ( .A(fifo_array[812]), .B(n4710), .Y(n1001) );
  INVX1 U266 ( .A(n1001), .Y(n149) );
  AND2X1 U268 ( .A(fifo_array[810]), .B(n4711), .Y(n999) );
  INVX1 U270 ( .A(n999), .Y(n150) );
  AND2X1 U272 ( .A(fifo_array[809]), .B(n4711), .Y(n998) );
  INVX1 U274 ( .A(n998), .Y(n151) );
  AND2X1 U276 ( .A(fifo_array[781]), .B(n4713), .Y(n969) );
  INVX1 U278 ( .A(n969), .Y(n152) );
  AND2X1 U280 ( .A(fifo_array[780]), .B(n4713), .Y(n968) );
  INVX1 U282 ( .A(n968), .Y(n153) );
  AND2X1 U284 ( .A(fifo_array[779]), .B(n4713), .Y(n967) );
  INVX1 U286 ( .A(n967), .Y(n1304) );
  AND2X1 U288 ( .A(fifo_array[778]), .B(n4712), .Y(n966) );
  INVX1 U290 ( .A(n966), .Y(n2464) );
  AND2X1 U292 ( .A(fifo_array[776]), .B(n4713), .Y(n964) );
  INVX1 U294 ( .A(n964), .Y(n2465) );
  AND2X1 U296 ( .A(fifo_array[775]), .B(n4713), .Y(n963) );
  INVX1 U298 ( .A(n963), .Y(n2466) );
  AND2X1 U300 ( .A(fifo_array[747]), .B(n4715), .Y(n934) );
  INVX1 U302 ( .A(n934), .Y(n2467) );
  AND2X1 U304 ( .A(fifo_array[746]), .B(n4715), .Y(n933) );
  INVX1 U306 ( .A(n933), .Y(n2468) );
  AND2X1 U308 ( .A(fifo_array[745]), .B(n4715), .Y(n932) );
  INVX1 U309 ( .A(n932), .Y(n2469) );
  AND2X1 U311 ( .A(fifo_array[744]), .B(n4714), .Y(n931) );
  INVX1 U313 ( .A(n931), .Y(n2470) );
  AND2X1 U315 ( .A(fifo_array[742]), .B(n4715), .Y(n929) );
  INVX1 U317 ( .A(n929), .Y(n2471) );
  AND2X1 U319 ( .A(fifo_array[741]), .B(n4715), .Y(n928) );
  INVX1 U321 ( .A(n928), .Y(n2472) );
  AND2X1 U323 ( .A(fifo_array[713]), .B(n4717), .Y(n899) );
  INVX1 U325 ( .A(n899), .Y(n2473) );
  AND2X1 U327 ( .A(fifo_array[712]), .B(n4717), .Y(n898) );
  INVX1 U329 ( .A(n898), .Y(n2474) );
  AND2X1 U331 ( .A(fifo_array[711]), .B(n4717), .Y(n897) );
  INVX1 U333 ( .A(n897), .Y(n2475) );
  AND2X1 U335 ( .A(fifo_array[710]), .B(n4716), .Y(n896) );
  INVX1 U337 ( .A(n896), .Y(n2476) );
  AND2X1 U339 ( .A(fifo_array[708]), .B(n4717), .Y(n894) );
  INVX1 U341 ( .A(n894), .Y(n2477) );
  AND2X1 U343 ( .A(fifo_array[707]), .B(n4717), .Y(n893) );
  INVX1 U345 ( .A(n893), .Y(n2478) );
  AND2X1 U347 ( .A(fifo_array[679]), .B(n4719), .Y(n864) );
  INVX1 U349 ( .A(n864), .Y(n2479) );
  AND2X1 U351 ( .A(fifo_array[678]), .B(n4719), .Y(n863) );
  INVX1 U353 ( .A(n863), .Y(n2480) );
  AND2X1 U355 ( .A(fifo_array[677]), .B(n4719), .Y(n862) );
  INVX1 U357 ( .A(n862), .Y(n2481) );
  AND2X1 U359 ( .A(fifo_array[676]), .B(n4718), .Y(n861) );
  INVX1 U361 ( .A(n861), .Y(n2482) );
  AND2X1 U363 ( .A(fifo_array[674]), .B(n4719), .Y(n859) );
  INVX1 U365 ( .A(n859), .Y(n2483) );
  AND2X1 U367 ( .A(fifo_array[673]), .B(n4719), .Y(n858) );
  INVX1 U369 ( .A(n858), .Y(n2484) );
  AND2X1 U371 ( .A(fifo_array[645]), .B(n4721), .Y(n829) );
  INVX1 U373 ( .A(n829), .Y(n2485) );
  AND2X1 U375 ( .A(fifo_array[644]), .B(n4721), .Y(n828) );
  INVX1 U377 ( .A(n828), .Y(n2486) );
  AND2X1 U378 ( .A(fifo_array[643]), .B(n4721), .Y(n827) );
  INVX1 U380 ( .A(n827), .Y(n2487) );
  AND2X1 U382 ( .A(fifo_array[642]), .B(n4720), .Y(n826) );
  INVX1 U384 ( .A(n826), .Y(n2488) );
  AND2X1 U386 ( .A(fifo_array[640]), .B(n4721), .Y(n824) );
  INVX1 U388 ( .A(n824), .Y(n2489) );
  AND2X1 U390 ( .A(fifo_array[639]), .B(n4721), .Y(n823) );
  INVX1 U392 ( .A(n823), .Y(n2490) );
  AND2X1 U394 ( .A(fifo_array[611]), .B(n4723), .Y(n794) );
  INVX1 U396 ( .A(n794), .Y(n2491) );
  AND2X1 U398 ( .A(fifo_array[610]), .B(n4723), .Y(n793) );
  INVX1 U400 ( .A(n793), .Y(n2492) );
  AND2X1 U402 ( .A(fifo_array[609]), .B(n4723), .Y(n792) );
  INVX1 U404 ( .A(n792), .Y(n2493) );
  AND2X1 U406 ( .A(fifo_array[608]), .B(n4722), .Y(n791) );
  INVX1 U408 ( .A(n791), .Y(n2494) );
  AND2X1 U410 ( .A(fifo_array[606]), .B(n4723), .Y(n789) );
  INVX1 U412 ( .A(n789), .Y(n2495) );
  AND2X1 U414 ( .A(fifo_array[605]), .B(n4723), .Y(n788) );
  INVX1 U416 ( .A(n788), .Y(n2496) );
  AND2X1 U418 ( .A(fifo_array[577]), .B(n4725), .Y(n758) );
  INVX1 U420 ( .A(n758), .Y(n2497) );
  AND2X1 U422 ( .A(fifo_array[576]), .B(n4725), .Y(n757) );
  INVX1 U424 ( .A(n757), .Y(n2498) );
  AND2X1 U426 ( .A(fifo_array[575]), .B(n4725), .Y(n756) );
  INVX1 U428 ( .A(n756), .Y(n2499) );
  AND2X1 U430 ( .A(fifo_array[574]), .B(n4724), .Y(n755) );
  INVX1 U432 ( .A(n755), .Y(n2500) );
  AND2X1 U434 ( .A(fifo_array[572]), .B(n4725), .Y(n753) );
  INVX1 U436 ( .A(n753), .Y(n2501) );
  AND2X1 U438 ( .A(fifo_array[571]), .B(n4725), .Y(n752) );
  INVX1 U440 ( .A(n752), .Y(n2502) );
  AND2X1 U442 ( .A(fifo_array[543]), .B(n4727), .Y(n723) );
  INVX1 U444 ( .A(n723), .Y(n2503) );
  AND2X1 U446 ( .A(fifo_array[542]), .B(n4727), .Y(n722) );
  INVX1 U447 ( .A(n722), .Y(n2504) );
  AND2X1 U449 ( .A(fifo_array[541]), .B(n4727), .Y(n721) );
  INVX1 U451 ( .A(n721), .Y(n2505) );
  AND2X1 U453 ( .A(fifo_array[540]), .B(n4726), .Y(n720) );
  INVX1 U455 ( .A(n720), .Y(n2506) );
  AND2X1 U457 ( .A(fifo_array[538]), .B(n4727), .Y(n718) );
  INVX1 U459 ( .A(n718), .Y(n2507) );
  AND2X1 U461 ( .A(fifo_array[537]), .B(n4727), .Y(n717) );
  INVX1 U463 ( .A(n717), .Y(n2508) );
  AND2X1 U465 ( .A(fifo_array[509]), .B(n4729), .Y(n688) );
  INVX1 U467 ( .A(n688), .Y(n2509) );
  AND2X1 U469 ( .A(fifo_array[508]), .B(n4729), .Y(n687) );
  INVX1 U471 ( .A(n687), .Y(n2510) );
  AND2X1 U473 ( .A(fifo_array[507]), .B(n4729), .Y(n686) );
  INVX1 U475 ( .A(n686), .Y(n2511) );
  AND2X1 U477 ( .A(fifo_array[506]), .B(n4728), .Y(n685) );
  INVX1 U479 ( .A(n685), .Y(n2512) );
  AND2X1 U481 ( .A(fifo_array[504]), .B(n4729), .Y(n683) );
  INVX1 U483 ( .A(n683), .Y(n2513) );
  AND2X1 U485 ( .A(fifo_array[503]), .B(n4729), .Y(n682) );
  INVX1 U487 ( .A(n682), .Y(n2514) );
  AND2X1 U489 ( .A(fifo_array[475]), .B(n4731), .Y(n653) );
  INVX1 U491 ( .A(n653), .Y(n2515) );
  AND2X1 U493 ( .A(fifo_array[474]), .B(n4731), .Y(n652) );
  INVX1 U495 ( .A(n652), .Y(n2516) );
  AND2X1 U497 ( .A(fifo_array[473]), .B(n4731), .Y(n651) );
  INVX1 U499 ( .A(n651), .Y(n2517) );
  AND2X1 U501 ( .A(fifo_array[472]), .B(n4730), .Y(n650) );
  INVX1 U503 ( .A(n650), .Y(n2518) );
  AND2X1 U505 ( .A(fifo_array[470]), .B(n4731), .Y(n648) );
  INVX1 U507 ( .A(n648), .Y(n2519) );
  AND2X1 U509 ( .A(fifo_array[469]), .B(n4731), .Y(n647) );
  INVX1 U511 ( .A(n647), .Y(n2520) );
  AND2X1 U513 ( .A(fifo_array[441]), .B(n4733), .Y(n618) );
  INVX1 U515 ( .A(n618), .Y(n2521) );
  AND2X1 U516 ( .A(fifo_array[440]), .B(n4733), .Y(n617) );
  INVX1 U518 ( .A(n617), .Y(n2522) );
  AND2X1 U520 ( .A(fifo_array[439]), .B(n4733), .Y(n616) );
  INVX1 U522 ( .A(n616), .Y(n2523) );
  AND2X1 U524 ( .A(fifo_array[438]), .B(n4732), .Y(n615) );
  INVX1 U526 ( .A(n615), .Y(n2524) );
  AND2X1 U528 ( .A(fifo_array[436]), .B(n4733), .Y(n613) );
  INVX1 U530 ( .A(n613), .Y(n2525) );
  AND2X1 U532 ( .A(fifo_array[435]), .B(n4733), .Y(n612) );
  INVX1 U534 ( .A(n612), .Y(n2526) );
  AND2X1 U536 ( .A(fifo_array[407]), .B(n4735), .Y(n583) );
  INVX1 U538 ( .A(n583), .Y(n2527) );
  AND2X1 U540 ( .A(fifo_array[406]), .B(n4735), .Y(n582) );
  INVX1 U542 ( .A(n582), .Y(n2528) );
  AND2X1 U544 ( .A(fifo_array[405]), .B(n4735), .Y(n581) );
  INVX1 U546 ( .A(n581), .Y(n2529) );
  AND2X1 U548 ( .A(fifo_array[404]), .B(n4734), .Y(n580) );
  INVX1 U550 ( .A(n580), .Y(n2530) );
  AND2X1 U552 ( .A(fifo_array[402]), .B(n4735), .Y(n578) );
  INVX1 U554 ( .A(n578), .Y(n2531) );
  AND2X1 U556 ( .A(fifo_array[401]), .B(n4735), .Y(n577) );
  INVX1 U558 ( .A(n577), .Y(n2532) );
  AND2X1 U560 ( .A(fifo_array[373]), .B(n4737), .Y(n548) );
  INVX1 U562 ( .A(n548), .Y(n2533) );
  AND2X1 U564 ( .A(fifo_array[372]), .B(n4737), .Y(n547) );
  INVX1 U566 ( .A(n547), .Y(n2534) );
  AND2X1 U568 ( .A(fifo_array[371]), .B(n4737), .Y(n546) );
  INVX1 U570 ( .A(n546), .Y(n2535) );
  AND2X1 U572 ( .A(fifo_array[370]), .B(n4736), .Y(n545) );
  INVX1 U574 ( .A(n545), .Y(n2536) );
  AND2X1 U576 ( .A(fifo_array[368]), .B(n4737), .Y(n543) );
  INVX1 U578 ( .A(n543), .Y(n2537) );
  AND2X1 U580 ( .A(fifo_array[367]), .B(n4737), .Y(n542) );
  INVX1 U582 ( .A(n542), .Y(n2538) );
  AND2X1 U584 ( .A(fifo_array[339]), .B(n4739), .Y(n513) );
  INVX1 U585 ( .A(n513), .Y(n2539) );
  AND2X1 U587 ( .A(fifo_array[338]), .B(n4739), .Y(n512) );
  INVX1 U589 ( .A(n512), .Y(n2540) );
  AND2X1 U591 ( .A(fifo_array[337]), .B(n4739), .Y(n511) );
  INVX1 U593 ( .A(n511), .Y(n2541) );
  AND2X1 U595 ( .A(fifo_array[336]), .B(n4738), .Y(n510) );
  INVX1 U597 ( .A(n510), .Y(n2542) );
  AND2X1 U599 ( .A(fifo_array[334]), .B(n4739), .Y(n508) );
  INVX1 U601 ( .A(n508), .Y(n2543) );
  AND2X1 U603 ( .A(fifo_array[333]), .B(n4739), .Y(n507) );
  INVX1 U605 ( .A(n507), .Y(n2544) );
  AND2X1 U607 ( .A(fifo_array[305]), .B(n4741), .Y(n477) );
  INVX1 U609 ( .A(n477), .Y(n2545) );
  AND2X1 U611 ( .A(fifo_array[304]), .B(n4741), .Y(n476) );
  INVX1 U613 ( .A(n476), .Y(n2546) );
  AND2X1 U615 ( .A(fifo_array[303]), .B(n4741), .Y(n475) );
  INVX1 U617 ( .A(n475), .Y(n2547) );
  AND2X1 U619 ( .A(fifo_array[302]), .B(n4740), .Y(n474) );
  INVX1 U621 ( .A(n474), .Y(n2548) );
  AND2X1 U623 ( .A(fifo_array[300]), .B(n4741), .Y(n472) );
  INVX1 U625 ( .A(n472), .Y(n2549) );
  AND2X1 U627 ( .A(fifo_array[299]), .B(n4741), .Y(n471) );
  INVX1 U629 ( .A(n471), .Y(n2550) );
  AND2X1 U631 ( .A(fifo_array[271]), .B(n4743), .Y(n441) );
  INVX1 U633 ( .A(n441), .Y(n2551) );
  AND2X1 U635 ( .A(fifo_array[270]), .B(n4743), .Y(n440) );
  INVX1 U637 ( .A(n440), .Y(n2552) );
  AND2X1 U639 ( .A(fifo_array[269]), .B(n4742), .Y(n439) );
  INVX1 U641 ( .A(n439), .Y(n2553) );
  AND2X1 U643 ( .A(fifo_array[268]), .B(n4743), .Y(n438) );
  INVX1 U645 ( .A(n438), .Y(n2554) );
  AND2X1 U647 ( .A(fifo_array[266]), .B(n4743), .Y(n436) );
  INVX1 U649 ( .A(n436), .Y(n2555) );
  AND2X1 U651 ( .A(fifo_array[265]), .B(n4743), .Y(n435) );
  INVX1 U653 ( .A(n435), .Y(n2556) );
  AND2X1 U654 ( .A(fifo_array[237]), .B(n4745), .Y(n405) );
  INVX1 U657 ( .A(n405), .Y(n2557) );
  AND2X1 U659 ( .A(fifo_array[236]), .B(n4745), .Y(n404) );
  INVX1 U661 ( .A(n404), .Y(n2558) );
  AND2X1 U663 ( .A(fifo_array[235]), .B(n4744), .Y(n403) );
  INVX1 U665 ( .A(n403), .Y(n2559) );
  AND2X1 U667 ( .A(fifo_array[234]), .B(n4745), .Y(n402) );
  INVX1 U669 ( .A(n402), .Y(n2560) );
  AND2X1 U671 ( .A(fifo_array[232]), .B(n4745), .Y(n400) );
  INVX1 U673 ( .A(n400), .Y(n2561) );
  AND2X1 U675 ( .A(fifo_array[231]), .B(n4745), .Y(n399) );
  INVX1 U677 ( .A(n399), .Y(n2562) );
  AND2X1 U679 ( .A(fifo_array[203]), .B(n4747), .Y(n369) );
  INVX1 U681 ( .A(n369), .Y(n2563) );
  AND2X1 U683 ( .A(fifo_array[202]), .B(n4747), .Y(n368) );
  INVX1 U685 ( .A(n368), .Y(n2564) );
  AND2X1 U687 ( .A(fifo_array[201]), .B(n4746), .Y(n367) );
  INVX1 U689 ( .A(n367), .Y(n2565) );
  AND2X1 U691 ( .A(fifo_array[200]), .B(n4747), .Y(n366) );
  INVX1 U693 ( .A(n366), .Y(n2566) );
  AND2X1 U695 ( .A(fifo_array[198]), .B(n4747), .Y(n364) );
  INVX1 U697 ( .A(n364), .Y(n2567) );
  AND2X1 U699 ( .A(fifo_array[197]), .B(n4747), .Y(n363) );
  INVX1 U701 ( .A(n363), .Y(n2568) );
  AND2X1 U703 ( .A(fifo_array[169]), .B(n4749), .Y(n333) );
  INVX1 U705 ( .A(n333), .Y(n2569) );
  AND2X1 U707 ( .A(fifo_array[168]), .B(n4749), .Y(n332) );
  INVX1 U709 ( .A(n332), .Y(n2570) );
  AND2X1 U711 ( .A(fifo_array[167]), .B(n4748), .Y(n331) );
  INVX1 U713 ( .A(n331), .Y(n2571) );
  AND2X1 U715 ( .A(fifo_array[166]), .B(n4749), .Y(n330) );
  INVX1 U717 ( .A(n330), .Y(n2572) );
  AND2X1 U719 ( .A(fifo_array[164]), .B(n4749), .Y(n328) );
  INVX1 U721 ( .A(n328), .Y(n2573) );
  AND2X1 U723 ( .A(fifo_array[163]), .B(n4749), .Y(n327) );
  INVX1 U724 ( .A(n327), .Y(n2574) );
  AND2X1 U726 ( .A(fifo_array[135]), .B(n4751), .Y(n297) );
  INVX1 U728 ( .A(n297), .Y(n2575) );
  AND2X1 U730 ( .A(fifo_array[134]), .B(n4751), .Y(n296) );
  INVX1 U732 ( .A(n296), .Y(n2576) );
  AND2X1 U734 ( .A(fifo_array[133]), .B(n4750), .Y(n295) );
  INVX1 U736 ( .A(n295), .Y(n2577) );
  AND2X1 U738 ( .A(fifo_array[132]), .B(n4751), .Y(n294) );
  INVX1 U740 ( .A(n294), .Y(n2578) );
  AND2X1 U742 ( .A(fifo_array[130]), .B(n4751), .Y(n292) );
  INVX1 U744 ( .A(n292), .Y(n2579) );
  AND2X1 U746 ( .A(fifo_array[129]), .B(n4751), .Y(n291) );
  INVX1 U748 ( .A(n291), .Y(n2580) );
  AND2X1 U750 ( .A(fifo_array[101]), .B(n4753), .Y(n261) );
  INVX1 U752 ( .A(n261), .Y(n2581) );
  AND2X1 U754 ( .A(fifo_array[100]), .B(n4753), .Y(n260) );
  INVX1 U756 ( .A(n260), .Y(n2582) );
  AND2X1 U758 ( .A(fifo_array[99]), .B(n4752), .Y(n259) );
  INVX1 U760 ( .A(n259), .Y(n2583) );
  AND2X1 U762 ( .A(fifo_array[98]), .B(n4753), .Y(n258) );
  INVX1 U764 ( .A(n258), .Y(n2584) );
  AND2X1 U766 ( .A(fifo_array[96]), .B(n4753), .Y(n256) );
  INVX1 U768 ( .A(n256), .Y(n2585) );
  AND2X1 U770 ( .A(fifo_array[95]), .B(n4753), .Y(n255) );
  INVX1 U772 ( .A(n255), .Y(n2586) );
  AND2X1 U774 ( .A(fifo_array[67]), .B(n4755), .Y(n225) );
  INVX1 U776 ( .A(n225), .Y(n2587) );
  AND2X1 U778 ( .A(fifo_array[66]), .B(n4755), .Y(n224) );
  INVX1 U780 ( .A(n224), .Y(n2588) );
  AND2X1 U782 ( .A(fifo_array[65]), .B(n4754), .Y(n223) );
  INVX1 U784 ( .A(n223), .Y(n2589) );
  AND2X1 U786 ( .A(fifo_array[64]), .B(n4755), .Y(n222) );
  INVX1 U788 ( .A(n222), .Y(n2590) );
  AND2X1 U790 ( .A(fifo_array[62]), .B(n4755), .Y(n220) );
  INVX1 U792 ( .A(n220), .Y(n2591) );
  AND2X1 U793 ( .A(fifo_array[61]), .B(n4755), .Y(n219) );
  INVX1 U795 ( .A(n219), .Y(n2592) );
  AND2X1 U797 ( .A(fifo_array[33]), .B(n4757), .Y(n188) );
  INVX1 U799 ( .A(n188), .Y(n2593) );
  AND2X1 U801 ( .A(fifo_array[32]), .B(n4757), .Y(n187) );
  INVX1 U803 ( .A(n187), .Y(n2594) );
  AND2X1 U805 ( .A(fifo_array[31]), .B(n4756), .Y(n186) );
  INVX1 U807 ( .A(n186), .Y(n2595) );
  AND2X1 U809 ( .A(fifo_array[30]), .B(n4757), .Y(n185) );
  INVX1 U811 ( .A(n185), .Y(n2596) );
  AND2X1 U813 ( .A(fifo_array[28]), .B(n4757), .Y(n183) );
  INVX1 U815 ( .A(n183), .Y(n2597) );
  AND2X1 U817 ( .A(fifo_array[27]), .B(n4757), .Y(n182) );
  INVX1 U819 ( .A(n182), .Y(n2598) );
  AND2X1 U821 ( .A(fifo_array[1076]), .B(n4694), .Y(n1274) );
  INVX1 U823 ( .A(n1274), .Y(n2599) );
  AND2X1 U825 ( .A(fifo_array[1065]), .B(n4695), .Y(n1263) );
  INVX1 U827 ( .A(n1263), .Y(n2600) );
  AND2X1 U829 ( .A(fifo_array[1049]), .B(n4697), .Y(n1246) );
  INVX1 U831 ( .A(n1246), .Y(n2601) );
  AND2X1 U833 ( .A(fifo_array[1032]), .B(n4697), .Y(n1229) );
  INVX1 U835 ( .A(n1229), .Y(n2602) );
  AND2X1 U837 ( .A(fifo_array[1009]), .B(n4699), .Y(n1205) );
  INVX1 U839 ( .A(n1205), .Y(n2603) );
  AND2X1 U841 ( .A(fifo_array[976]), .B(n4701), .Y(n1171) );
  INVX1 U843 ( .A(n1171), .Y(n2604) );
  AND2X1 U845 ( .A(fifo_array[943]), .B(n4703), .Y(n1137) );
  INVX1 U847 ( .A(n1137), .Y(n2605) );
  AND2X1 U849 ( .A(fifo_array[910]), .B(n4705), .Y(n1103) );
  INVX1 U851 ( .A(n1103), .Y(n2606) );
  AND2X1 U853 ( .A(fifo_array[865]), .B(n4707), .Y(n1057) );
  INVX1 U855 ( .A(n1057), .Y(n2607) );
  AND2X1 U857 ( .A(fifo_array[853]), .B(n4707), .Y(n1045) );
  INVX1 U859 ( .A(n1045), .Y(n2608) );
  AND2X1 U861 ( .A(fifo_array[832]), .B(n4709), .Y(n1022) );
  INVX1 U862 ( .A(n1022), .Y(n2609) );
  AND2X1 U864 ( .A(fifo_array[820]), .B(n4709), .Y(n1010) );
  INVX1 U866 ( .A(n1010), .Y(n2610) );
  AND2X1 U868 ( .A(fifo_array[799]), .B(n4711), .Y(n988) );
  INVX1 U870 ( .A(n988), .Y(n2611) );
  AND2X1 U872 ( .A(fifo_array[787]), .B(n4710), .Y(n976) );
  INVX1 U874 ( .A(n976), .Y(n2612) );
  AND2X1 U876 ( .A(fifo_array[766]), .B(n4713), .Y(n954) );
  INVX1 U878 ( .A(n954), .Y(n2613) );
  AND2X1 U880 ( .A(fifo_array[754]), .B(n4712), .Y(n942) );
  INVX1 U882 ( .A(n942), .Y(n2614) );
  AND2X1 U884 ( .A(fifo_array[733]), .B(n4715), .Y(n920) );
  INVX1 U886 ( .A(n920), .Y(n2615) );
  AND2X1 U888 ( .A(fifo_array[721]), .B(n4714), .Y(n908) );
  INVX1 U890 ( .A(n908), .Y(n2616) );
  AND2X1 U892 ( .A(fifo_array[700]), .B(n4716), .Y(n886) );
  INVX1 U894 ( .A(n886), .Y(n2617) );
  AND2X1 U896 ( .A(fifo_array[688]), .B(n4716), .Y(n874) );
  INVX1 U898 ( .A(n874), .Y(n2618) );
  AND2X1 U900 ( .A(fifo_array[667]), .B(n4718), .Y(n852) );
  INVX1 U902 ( .A(n852), .Y(n2619) );
  AND2X1 U904 ( .A(fifo_array[656]), .B(n4719), .Y(n841) );
  INVX1 U906 ( .A(n841), .Y(n2620) );
  AND2X1 U908 ( .A(fifo_array[634]), .B(n4720), .Y(n818) );
  INVX1 U910 ( .A(n818), .Y(n2621) );
  AND2X1 U912 ( .A(fifo_array[623]), .B(n4721), .Y(n807) );
  INVX1 U914 ( .A(n807), .Y(n2622) );
  AND2X1 U916 ( .A(fifo_array[607]), .B(n4722), .Y(n790) );
  INVX1 U918 ( .A(n790), .Y(n2623) );
  AND2X1 U920 ( .A(fifo_array[590]), .B(n4723), .Y(n773) );
  INVX1 U922 ( .A(n773), .Y(n2624) );
  AND2X1 U924 ( .A(fifo_array[567]), .B(n4725), .Y(n748) );
  INVX1 U926 ( .A(n748), .Y(n2625) );
  AND2X1 U928 ( .A(fifo_array[534]), .B(n4727), .Y(n714) );
  INVX1 U930 ( .A(n714), .Y(n2626) );
  AND2X1 U931 ( .A(fifo_array[501]), .B(n4729), .Y(n680) );
  INVX1 U933 ( .A(n680), .Y(n2627) );
  AND2X1 U935 ( .A(fifo_array[468]), .B(n4731), .Y(n646) );
  INVX1 U937 ( .A(n646), .Y(n2628) );
  AND2X1 U939 ( .A(fifo_array[423]), .B(n4733), .Y(n600) );
  INVX1 U941 ( .A(n600), .Y(n2629) );
  AND2X1 U943 ( .A(fifo_array[411]), .B(n4732), .Y(n588) );
  INVX1 U945 ( .A(n588), .Y(n2630) );
  AND2X1 U947 ( .A(fifo_array[390]), .B(n4735), .Y(n566) );
  INVX1 U949 ( .A(n566), .Y(n2631) );
  AND2X1 U951 ( .A(fifo_array[378]), .B(n4734), .Y(n554) );
  INVX1 U953 ( .A(n554), .Y(n2632) );
  AND2X1 U955 ( .A(fifo_array[357]), .B(n4737), .Y(n532) );
  INVX1 U957 ( .A(n532), .Y(n2633) );
  AND2X1 U959 ( .A(fifo_array[345]), .B(n4736), .Y(n520) );
  INVX1 U961 ( .A(n520), .Y(n2634) );
  AND2X1 U963 ( .A(fifo_array[324]), .B(n4739), .Y(n498) );
  INVX1 U965 ( .A(n498), .Y(n2635) );
  AND2X1 U967 ( .A(fifo_array[312]), .B(n4738), .Y(n486) );
  INVX1 U969 ( .A(n486), .Y(n2636) );
  AND2X1 U971 ( .A(fifo_array[291]), .B(n4741), .Y(n463) );
  INVX1 U973 ( .A(n463), .Y(n2637) );
  AND2X1 U975 ( .A(fifo_array[279]), .B(n4740), .Y(n451) );
  INVX1 U977 ( .A(n451), .Y(n2638) );
  AND2X1 U979 ( .A(fifo_array[258]), .B(n4742), .Y(n428) );
  INVX1 U981 ( .A(n428), .Y(n2639) );
  AND2X1 U983 ( .A(fifo_array[246]), .B(n4743), .Y(n416) );
  INVX1 U985 ( .A(n416), .Y(n2640) );
  AND2X1 U987 ( .A(fifo_array[225]), .B(n4744), .Y(n393) );
  INVX1 U989 ( .A(n393), .Y(n2641) );
  AND2X1 U991 ( .A(fifo_array[214]), .B(n4745), .Y(n382) );
  INVX1 U993 ( .A(n382), .Y(n2642) );
  AND2X1 U995 ( .A(fifo_array[192]), .B(n4746), .Y(n358) );
  INVX1 U997 ( .A(n358), .Y(n2643) );
  AND2X1 U999 ( .A(fifo_array[181]), .B(n4747), .Y(n347) );
  INVX1 U1000 ( .A(n347), .Y(n2644) );
  AND2X1 U1002 ( .A(fifo_array[165]), .B(n4749), .Y(n329) );
  INVX1 U1004 ( .A(n329), .Y(n2645) );
  AND2X1 U1006 ( .A(fifo_array[148]), .B(n4749), .Y(n312) );
  INVX1 U1008 ( .A(n312), .Y(n2646) );
  AND2X1 U1010 ( .A(fifo_array[125]), .B(n4751), .Y(n287) );
  INVX1 U1012 ( .A(n287), .Y(n2647) );
  AND2X1 U1014 ( .A(fifo_array[92]), .B(n4753), .Y(n252) );
  INVX1 U1016 ( .A(n252), .Y(n2648) );
  AND2X1 U1018 ( .A(fifo_array[59]), .B(n4755), .Y(n217) );
  INVX1 U1020 ( .A(n217), .Y(n2649) );
  AND2X1 U1022 ( .A(fifo_array[26]), .B(n4757), .Y(n181) );
  INVX1 U1024 ( .A(n181), .Y(n2650) );
  AND2X1 U1026 ( .A(fifo_array[1083]), .B(n4695), .Y(n1281) );
  INVX1 U1028 ( .A(n1281), .Y(n2651) );
  AND2X1 U1030 ( .A(fifo_array[1066]), .B(n4695), .Y(n1264) );
  INVX1 U1032 ( .A(n1264), .Y(n2652) );
  AND2X1 U1034 ( .A(fifo_array[1042]), .B(n4696), .Y(n1239) );
  INVX1 U1036 ( .A(n1239), .Y(n2653) );
  AND2X1 U1038 ( .A(fifo_array[1031]), .B(n4697), .Y(n1228) );
  INVX1 U1040 ( .A(n1228), .Y(n2654) );
  AND2X1 U1042 ( .A(fifo_array[1010]), .B(n4699), .Y(n1206) );
  INVX1 U1044 ( .A(n1206), .Y(n2655) );
  AND2X1 U1046 ( .A(fifo_array[975]), .B(n4701), .Y(n1170) );
  INVX1 U1048 ( .A(n1170), .Y(n2656) );
  AND2X1 U1050 ( .A(fifo_array[944]), .B(n4703), .Y(n1138) );
  INVX1 U1052 ( .A(n1138), .Y(n2657) );
  AND2X1 U1054 ( .A(fifo_array[909]), .B(n4705), .Y(n1102) );
  INVX1 U1056 ( .A(n1102), .Y(n2658) );
  AND2X1 U1058 ( .A(fifo_array[864]), .B(n4707), .Y(n1056) );
  INVX1 U1060 ( .A(n1056), .Y(n2659) );
  AND2X1 U1062 ( .A(fifo_array[852]), .B(n4707), .Y(n1044) );
  INVX1 U1064 ( .A(n1044), .Y(n2660) );
  AND2X1 U1066 ( .A(fifo_array[833]), .B(n4709), .Y(n1023) );
  INVX1 U1068 ( .A(n1023), .Y(n2661) );
  AND2X1 U1069 ( .A(fifo_array[821]), .B(n4709), .Y(n1011) );
  INVX1 U1071 ( .A(n1011), .Y(n2662) );
  AND2X1 U1073 ( .A(fifo_array[798]), .B(n4711), .Y(n987) );
  INVX1 U1075 ( .A(n987), .Y(n2663) );
  AND2X1 U1077 ( .A(fifo_array[786]), .B(n4711), .Y(n975) );
  INVX1 U1079 ( .A(n975), .Y(n2664) );
  AND2X1 U1081 ( .A(fifo_array[767]), .B(n4713), .Y(n955) );
  INVX1 U1083 ( .A(n955), .Y(n2665) );
  AND2X1 U1085 ( .A(fifo_array[755]), .B(n4713), .Y(n943) );
  INVX1 U1087 ( .A(n943), .Y(n2666) );
  AND2X1 U1089 ( .A(fifo_array[732]), .B(n4715), .Y(n919) );
  INVX1 U1091 ( .A(n919), .Y(n2667) );
  AND2X1 U1093 ( .A(fifo_array[720]), .B(n4715), .Y(n907) );
  INVX1 U1095 ( .A(n907), .Y(n2668) );
  AND2X1 U1097 ( .A(fifo_array[701]), .B(n4716), .Y(n887) );
  INVX1 U1099 ( .A(n887), .Y(n2669) );
  AND2X1 U1101 ( .A(fifo_array[690]), .B(n4717), .Y(n876) );
  INVX1 U1103 ( .A(n876), .Y(n2670) );
  AND2X1 U1105 ( .A(fifo_array[666]), .B(n4718), .Y(n851) );
  INVX1 U1107 ( .A(n851), .Y(n2671) );
  AND2X1 U1109 ( .A(fifo_array[654]), .B(n4718), .Y(n839) );
  INVX1 U1111 ( .A(n839), .Y(n2672) );
  AND2X1 U1113 ( .A(fifo_array[641]), .B(n4720), .Y(n825) );
  INVX1 U1115 ( .A(n825), .Y(n2673) );
  AND2X1 U1117 ( .A(fifo_array[624]), .B(n4721), .Y(n808) );
  INVX1 U1119 ( .A(n808), .Y(n2674) );
  AND2X1 U1121 ( .A(fifo_array[600]), .B(n4722), .Y(n783) );
  INVX1 U1123 ( .A(n783), .Y(n2675) );
  AND2X1 U1125 ( .A(fifo_array[589]), .B(n4723), .Y(n772) );
  INVX1 U1127 ( .A(n772), .Y(n2676) );
  AND2X1 U1129 ( .A(fifo_array[568]), .B(n4725), .Y(n749) );
  INVX1 U1131 ( .A(n749), .Y(n2677) );
  AND2X1 U1133 ( .A(fifo_array[533]), .B(n4727), .Y(n713) );
  INVX1 U1135 ( .A(n713), .Y(n2678) );
  AND2X1 U1137 ( .A(fifo_array[502]), .B(n4729), .Y(n681) );
  INVX1 U1138 ( .A(n681), .Y(n2679) );
  AND2X1 U1140 ( .A(fifo_array[467]), .B(n4731), .Y(n645) );
  INVX1 U1142 ( .A(n645), .Y(n2680) );
  AND2X1 U1144 ( .A(fifo_array[422]), .B(n4733), .Y(n599) );
  INVX1 U1146 ( .A(n599), .Y(n2681) );
  AND2X1 U1148 ( .A(fifo_array[410]), .B(n4733), .Y(n587) );
  INVX1 U1150 ( .A(n587), .Y(n2682) );
  AND2X1 U1152 ( .A(fifo_array[391]), .B(n4735), .Y(n567) );
  INVX1 U1154 ( .A(n567), .Y(n2683) );
  AND2X1 U1156 ( .A(fifo_array[379]), .B(n4735), .Y(n555) );
  INVX1 U1158 ( .A(n555), .Y(n2684) );
  AND2X1 U1160 ( .A(fifo_array[356]), .B(n4737), .Y(n531) );
  INVX1 U1162 ( .A(n531), .Y(n2685) );
  AND2X1 U1164 ( .A(fifo_array[344]), .B(n4737), .Y(n519) );
  INVX1 U1166 ( .A(n519), .Y(n2686) );
  AND2X1 U1168 ( .A(fifo_array[325]), .B(n4739), .Y(n499) );
  INVX1 U1170 ( .A(n499), .Y(n2687) );
  AND2X1 U1172 ( .A(fifo_array[313]), .B(n4739), .Y(n487) );
  INVX1 U1174 ( .A(n487), .Y(n2688) );
  AND2X1 U1176 ( .A(fifo_array[290]), .B(n4741), .Y(n462) );
  INVX1 U1178 ( .A(n462), .Y(n2689) );
  AND2X1 U1180 ( .A(fifo_array[278]), .B(n4741), .Y(n450) );
  INVX1 U1182 ( .A(n450), .Y(n2690) );
  AND2X1 U1184 ( .A(fifo_array[259]), .B(n4743), .Y(n429) );
  INVX1 U1186 ( .A(n429), .Y(n2691) );
  AND2X1 U1188 ( .A(fifo_array[248]), .B(n4743), .Y(n418) );
  INVX1 U1190 ( .A(n418), .Y(n2692) );
  AND2X1 U1192 ( .A(fifo_array[224]), .B(n4745), .Y(n392) );
  INVX1 U1194 ( .A(n392), .Y(n2693) );
  AND2X1 U1196 ( .A(fifo_array[212]), .B(n4745), .Y(n380) );
  INVX1 U1198 ( .A(n380), .Y(n2694) );
  AND2X1 U1200 ( .A(fifo_array[199]), .B(n4747), .Y(n365) );
  INVX1 U1202 ( .A(n365), .Y(n2695) );
  AND2X1 U1204 ( .A(fifo_array[182]), .B(n4747), .Y(n348) );
  INVX1 U1206 ( .A(n348), .Y(n2696) );
  AND2X1 U1207 ( .A(fifo_array[158]), .B(n4748), .Y(n322) );
  INVX1 U1210 ( .A(n322), .Y(n2697) );
  AND2X1 U1212 ( .A(fifo_array[147]), .B(n4749), .Y(n311) );
  INVX1 U1214 ( .A(n311), .Y(n2698) );
  AND2X1 U1216 ( .A(fifo_array[126]), .B(n4751), .Y(n288) );
  INVX1 U1218 ( .A(n288), .Y(n2699) );
  AND2X1 U1220 ( .A(fifo_array[91]), .B(n4753), .Y(n251) );
  INVX1 U1222 ( .A(n251), .Y(n2700) );
  AND2X1 U1224 ( .A(fifo_array[60]), .B(n4755), .Y(n218) );
  INVX1 U1226 ( .A(n218), .Y(n2701) );
  AND2X1 U1228 ( .A(fifo_array[25]), .B(n4757), .Y(n180) );
  INVX1 U1230 ( .A(n180), .Y(n2702) );
  AND2X1 U1232 ( .A(fifo_array[1074]), .B(n4694), .Y(n1272) );
  INVX1 U1234 ( .A(n1272), .Y(n2703) );
  AND2X1 U1236 ( .A(fifo_array[1062]), .B(n4695), .Y(n1260) );
  INVX1 U1238 ( .A(n1260), .Y(n2704) );
  AND2X1 U1240 ( .A(fifo_array[1041]), .B(n4696), .Y(n1238) );
  INVX1 U1242 ( .A(n1238), .Y(n2705) );
  AND2X1 U1244 ( .A(fifo_array[1030]), .B(n4697), .Y(n1227) );
  INVX1 U1246 ( .A(n1227), .Y(n2706) );
  AND2X1 U1248 ( .A(fifo_array[1011]), .B(n4699), .Y(n1207) );
  INVX1 U1250 ( .A(n1207), .Y(n2707) );
  AND2X1 U1252 ( .A(fifo_array[978]), .B(n4701), .Y(n1173) );
  INVX1 U1254 ( .A(n1173), .Y(n2708) );
  AND2X1 U1256 ( .A(fifo_array[941]), .B(n4703), .Y(n1135) );
  INVX1 U1258 ( .A(n1135), .Y(n2709) );
  AND2X1 U1260 ( .A(fifo_array[908]), .B(n4705), .Y(n1101) );
  INVX1 U1262 ( .A(n1101), .Y(n2710) );
  AND2X1 U1264 ( .A(fifo_array[863]), .B(n4707), .Y(n1055) );
  INVX1 U1266 ( .A(n1055), .Y(n2711) );
  AND2X1 U1268 ( .A(fifo_array[851]), .B(n4707), .Y(n1043) );
  INVX1 U1270 ( .A(n1043), .Y(n2712) );
  AND2X1 U1272 ( .A(fifo_array[834]), .B(n4709), .Y(n1024) );
  INVX1 U1274 ( .A(n1024), .Y(n2713) );
  AND2X1 U1276 ( .A(fifo_array[822]), .B(n4709), .Y(n1012) );
  INVX1 U1277 ( .A(n1012), .Y(n2714) );
  AND2X1 U1279 ( .A(fifo_array[801]), .B(n4711), .Y(n990) );
  INVX1 U1281 ( .A(n990), .Y(n2715) );
  AND2X1 U1283 ( .A(fifo_array[789]), .B(n4711), .Y(n978) );
  INVX1 U1285 ( .A(n978), .Y(n2716) );
  AND2X1 U1287 ( .A(fifo_array[764]), .B(n4713), .Y(n952) );
  INVX1 U1289 ( .A(n952), .Y(n2717) );
  AND2X1 U1291 ( .A(fifo_array[752]), .B(n4713), .Y(n940) );
  INVX1 U1293 ( .A(n940), .Y(n2718) );
  AND2X1 U1295 ( .A(fifo_array[731]), .B(n4715), .Y(n918) );
  INVX1 U1297 ( .A(n918), .Y(n2719) );
  AND2X1 U1299 ( .A(fifo_array[719]), .B(n4715), .Y(n906) );
  INVX1 U1301 ( .A(n906), .Y(n2720) );
  AND2X1 U1303 ( .A(fifo_array[702]), .B(n4716), .Y(n888) );
  INVX1 U1305 ( .A(n888), .Y(n2721) );
  AND2X1 U1307 ( .A(fifo_array[691]), .B(n4717), .Y(n877) );
  INVX1 U1309 ( .A(n877), .Y(n2722) );
  AND2X1 U1311 ( .A(fifo_array[675]), .B(n4719), .Y(n860) );
  INVX1 U1313 ( .A(n860), .Y(n2723) );
  AND2X1 U1315 ( .A(fifo_array[658]), .B(n4719), .Y(n843) );
  INVX1 U1317 ( .A(n843), .Y(n2724) );
  AND2X1 U1319 ( .A(fifo_array[632]), .B(n4720), .Y(n816) );
  INVX1 U1321 ( .A(n816), .Y(n2725) );
  AND2X1 U1323 ( .A(fifo_array[620]), .B(n4721), .Y(n804) );
  INVX1 U1325 ( .A(n804), .Y(n2726) );
  AND2X1 U1327 ( .A(fifo_array[599]), .B(n4722), .Y(n782) );
  INVX1 U1329 ( .A(n782), .Y(n2727) );
  AND2X1 U1331 ( .A(fifo_array[588]), .B(n4723), .Y(n771) );
  INVX1 U1333 ( .A(n771), .Y(n2728) );
  AND2X1 U1335 ( .A(fifo_array[569]), .B(n4725), .Y(n750) );
  INVX1 U1337 ( .A(n750), .Y(n2729) );
  AND2X1 U1339 ( .A(fifo_array[536]), .B(n4727), .Y(n716) );
  INVX1 U1341 ( .A(n716), .Y(n2730) );
  AND2X1 U1343 ( .A(fifo_array[499]), .B(n4729), .Y(n678) );
  INVX1 U1345 ( .A(n678), .Y(n2731) );
  AND2X1 U1346 ( .A(fifo_array[466]), .B(n4731), .Y(n644) );
  INVX1 U1348 ( .A(n644), .Y(n2732) );
  AND2X1 U1350 ( .A(fifo_array[421]), .B(n4733), .Y(n598) );
  INVX1 U1352 ( .A(n598), .Y(n2733) );
  AND2X1 U1354 ( .A(fifo_array[409]), .B(n4733), .Y(n586) );
  INVX1 U1356 ( .A(n586), .Y(n2734) );
  AND2X1 U1358 ( .A(fifo_array[392]), .B(n4735), .Y(n568) );
  INVX1 U1360 ( .A(n568), .Y(n2735) );
  AND2X1 U1362 ( .A(fifo_array[380]), .B(n4735), .Y(n556) );
  INVX1 U1364 ( .A(n556), .Y(n2736) );
  AND2X1 U1366 ( .A(fifo_array[359]), .B(n4737), .Y(n534) );
  INVX1 U1368 ( .A(n534), .Y(n2737) );
  AND2X1 U1370 ( .A(fifo_array[347]), .B(n4737), .Y(n522) );
  INVX1 U1372 ( .A(n522), .Y(n2738) );
  AND2X1 U1374 ( .A(fifo_array[322]), .B(n4739), .Y(n496) );
  INVX1 U1376 ( .A(n496), .Y(n2739) );
  AND2X1 U1378 ( .A(fifo_array[310]), .B(n4739), .Y(n484) );
  INVX1 U1380 ( .A(n484), .Y(n2740) );
  AND2X1 U1382 ( .A(fifo_array[289]), .B(n4741), .Y(n461) );
  INVX1 U1384 ( .A(n461), .Y(n2741) );
  AND2X1 U1386 ( .A(fifo_array[277]), .B(n4741), .Y(n449) );
  INVX1 U1388 ( .A(n449), .Y(n2742) );
  AND2X1 U1390 ( .A(fifo_array[260]), .B(n4743), .Y(n430) );
  INVX1 U1392 ( .A(n430), .Y(n2743) );
  AND2X1 U1394 ( .A(fifo_array[249]), .B(n4743), .Y(n419) );
  INVX1 U1396 ( .A(n419), .Y(n2744) );
  AND2X1 U1398 ( .A(fifo_array[233]), .B(n4745), .Y(n401) );
  INVX1 U1400 ( .A(n401), .Y(n2745) );
  AND2X1 U1402 ( .A(fifo_array[216]), .B(n4745), .Y(n384) );
  INVX1 U1404 ( .A(n384), .Y(n2746) );
  AND2X1 U1406 ( .A(fifo_array[190]), .B(n4747), .Y(n356) );
  INVX1 U1408 ( .A(n356), .Y(n2747) );
  AND2X1 U1410 ( .A(fifo_array[178]), .B(n4747), .Y(n344) );
  INVX1 U1412 ( .A(n344), .Y(n2748) );
  AND2X1 U1414 ( .A(fifo_array[157]), .B(n4749), .Y(n321) );
  INVX1 U1415 ( .A(n321), .Y(n2749) );
  AND2X1 U1417 ( .A(fifo_array[146]), .B(n4749), .Y(n310) );
  INVX1 U1419 ( .A(n310), .Y(n2750) );
  AND2X1 U1421 ( .A(fifo_array[127]), .B(n4751), .Y(n289) );
  INVX1 U1423 ( .A(n289), .Y(n2751) );
  AND2X1 U1425 ( .A(fifo_array[94]), .B(n4753), .Y(n254) );
  INVX1 U1427 ( .A(n254), .Y(n2752) );
  AND2X1 U1429 ( .A(fifo_array[57]), .B(n4755), .Y(n215) );
  INVX1 U1431 ( .A(n215), .Y(n2753) );
  AND2X1 U1433 ( .A(fifo_array[24]), .B(n4757), .Y(n179) );
  INVX1 U1435 ( .A(n179), .Y(n2754) );
  AND2X1 U1437 ( .A(fifo_array[1075]), .B(n4694), .Y(n1273) );
  INVX1 U1439 ( .A(n1273), .Y(n2755) );
  AND2X1 U1441 ( .A(fifo_array[1064]), .B(n4695), .Y(n1262) );
  INVX1 U1443 ( .A(n1262), .Y(n2756) );
  AND2X1 U1445 ( .A(fifo_array[1040]), .B(n4696), .Y(n1237) );
  INVX1 U1447 ( .A(n1237), .Y(n2757) );
  AND2X1 U1449 ( .A(fifo_array[1028]), .B(n4697), .Y(n1225) );
  INVX1 U1451 ( .A(n1225), .Y(n2758) );
  AND2X1 U1453 ( .A(fifo_array[1012]), .B(n4699), .Y(n1208) );
  INVX1 U1455 ( .A(n1208), .Y(n2759) );
  AND2X1 U1457 ( .A(fifo_array[977]), .B(n4701), .Y(n1172) );
  INVX1 U1459 ( .A(n1172), .Y(n2760) );
  AND2X1 U1461 ( .A(fifo_array[942]), .B(n4703), .Y(n1136) );
  INVX1 U1463 ( .A(n1136), .Y(n2761) );
  AND2X1 U1465 ( .A(fifo_array[907]), .B(n4705), .Y(n1100) );
  INVX1 U1467 ( .A(n1100), .Y(n2762) );
  AND2X1 U1469 ( .A(fifo_array[859]), .B(n4707), .Y(n1051) );
  INVX1 U1471 ( .A(n1051), .Y(n2763) );
  AND2X1 U1473 ( .A(fifo_array[850]), .B(n4706), .Y(n1042) );
  INVX1 U1475 ( .A(n1042), .Y(n2764) );
  AND2X1 U1477 ( .A(fifo_array[835]), .B(n4709), .Y(n1025) );
  INVX1 U1479 ( .A(n1025), .Y(n2765) );
  AND2X1 U1481 ( .A(fifo_array[823]), .B(n4708), .Y(n1013) );
  INVX1 U1483 ( .A(n1013), .Y(n2766) );
  AND2X1 U1484 ( .A(fifo_array[800]), .B(n4711), .Y(n989) );
  INVX1 U1486 ( .A(n989), .Y(n2767) );
  AND2X1 U1488 ( .A(fifo_array[788]), .B(n4710), .Y(n977) );
  INVX1 U1490 ( .A(n977), .Y(n2768) );
  AND2X1 U1492 ( .A(fifo_array[765]), .B(n4713), .Y(n953) );
  INVX1 U1494 ( .A(n953), .Y(n2769) );
  AND2X1 U1496 ( .A(fifo_array[753]), .B(n4712), .Y(n941) );
  INVX1 U1498 ( .A(n941), .Y(n2770) );
  AND2X1 U1500 ( .A(fifo_array[730]), .B(n4715), .Y(n917) );
  INVX1 U1502 ( .A(n917), .Y(n2771) );
  AND2X1 U1504 ( .A(fifo_array[718]), .B(n4714), .Y(n905) );
  INVX1 U1506 ( .A(n905), .Y(n2772) );
  AND2X1 U1508 ( .A(fifo_array[709]), .B(n4717), .Y(n895) );
  INVX1 U1510 ( .A(n895), .Y(n2773) );
  AND2X1 U1512 ( .A(fifo_array[692]), .B(n4717), .Y(n878) );
  INVX1 U1514 ( .A(n878), .Y(n2774) );
  AND2X1 U1516 ( .A(fifo_array[668]), .B(n4718), .Y(n853) );
  INVX1 U1518 ( .A(n853), .Y(n2775) );
  AND2X1 U1520 ( .A(fifo_array[657]), .B(n4719), .Y(n842) );
  INVX1 U1522 ( .A(n842), .Y(n2776) );
  AND2X1 U1524 ( .A(fifo_array[633]), .B(n4720), .Y(n817) );
  INVX1 U1526 ( .A(n817), .Y(n2777) );
  AND2X1 U1528 ( .A(fifo_array[622]), .B(n4721), .Y(n806) );
  INVX1 U1530 ( .A(n806), .Y(n2778) );
  AND2X1 U1532 ( .A(fifo_array[598]), .B(n4722), .Y(n781) );
  INVX1 U1534 ( .A(n781), .Y(n2779) );
  AND2X1 U1536 ( .A(fifo_array[586]), .B(n4723), .Y(n769) );
  INVX1 U1538 ( .A(n769), .Y(n2780) );
  AND2X1 U1540 ( .A(fifo_array[570]), .B(n4725), .Y(n751) );
  INVX1 U1542 ( .A(n751), .Y(n2781) );
  AND2X1 U1544 ( .A(fifo_array[535]), .B(n4727), .Y(n715) );
  INVX1 U1546 ( .A(n715), .Y(n2782) );
  AND2X1 U1548 ( .A(fifo_array[500]), .B(n4729), .Y(n679) );
  INVX1 U1550 ( .A(n679), .Y(n2783) );
  AND2X1 U1552 ( .A(fifo_array[465]), .B(n4731), .Y(n643) );
  INVX1 U1553 ( .A(n643), .Y(n2784) );
  AND2X1 U1555 ( .A(fifo_array[417]), .B(n4733), .Y(n594) );
  INVX1 U1557 ( .A(n594), .Y(n2785) );
  AND2X1 U1559 ( .A(fifo_array[408]), .B(n4732), .Y(n585) );
  INVX1 U1561 ( .A(n585), .Y(n2786) );
  AND2X1 U1563 ( .A(fifo_array[393]), .B(n4735), .Y(n569) );
  INVX1 U1565 ( .A(n569), .Y(n2787) );
  AND2X1 U1567 ( .A(fifo_array[381]), .B(n4734), .Y(n557) );
  INVX1 U1569 ( .A(n557), .Y(n2788) );
  AND2X1 U1571 ( .A(fifo_array[358]), .B(n4737), .Y(n533) );
  INVX1 U1573 ( .A(n533), .Y(n2789) );
  AND2X1 U1575 ( .A(fifo_array[346]), .B(n4736), .Y(n521) );
  INVX1 U1577 ( .A(n521), .Y(n2790) );
  AND2X1 U1579 ( .A(fifo_array[323]), .B(n4739), .Y(n497) );
  INVX1 U1581 ( .A(n497), .Y(n2791) );
  AND2X1 U1583 ( .A(fifo_array[311]), .B(n4738), .Y(n485) );
  INVX1 U1585 ( .A(n485), .Y(n2792) );
  AND2X1 U1587 ( .A(fifo_array[288]), .B(n4741), .Y(n460) );
  INVX1 U1589 ( .A(n460), .Y(n2793) );
  AND2X1 U1591 ( .A(fifo_array[276]), .B(n4740), .Y(n448) );
  INVX1 U1593 ( .A(n448), .Y(n2794) );
  AND2X1 U1595 ( .A(fifo_array[267]), .B(n4743), .Y(n437) );
  INVX1 U1597 ( .A(n437), .Y(n2795) );
  AND2X1 U1599 ( .A(fifo_array[250]), .B(n4743), .Y(n420) );
  INVX1 U1601 ( .A(n420), .Y(n2796) );
  AND2X1 U1603 ( .A(fifo_array[226]), .B(n4745), .Y(n394) );
  INVX1 U1605 ( .A(n394), .Y(n2797) );
  AND2X1 U1607 ( .A(fifo_array[215]), .B(n4745), .Y(n383) );
  INVX1 U1609 ( .A(n383), .Y(n2798) );
  AND2X1 U1611 ( .A(fifo_array[191]), .B(n4747), .Y(n357) );
  INVX1 U1613 ( .A(n357), .Y(n2799) );
  AND2X1 U1615 ( .A(fifo_array[180]), .B(n4747), .Y(n346) );
  INVX1 U1617 ( .A(n346), .Y(n2800) );
  AND2X1 U1619 ( .A(fifo_array[156]), .B(n4749), .Y(n320) );
  INVX1 U1621 ( .A(n320), .Y(n2801) );
  AND2X1 U1622 ( .A(fifo_array[144]), .B(n4749), .Y(n308) );
  INVX1 U1624 ( .A(n308), .Y(n2802) );
  AND2X1 U1626 ( .A(fifo_array[128]), .B(n4751), .Y(n290) );
  INVX1 U1628 ( .A(n290), .Y(n2803) );
  AND2X1 U1630 ( .A(fifo_array[93]), .B(n4753), .Y(n253) );
  INVX1 U1632 ( .A(n253), .Y(n2804) );
  AND2X1 U1634 ( .A(fifo_array[58]), .B(n4755), .Y(n216) );
  INVX1 U1636 ( .A(n216), .Y(n2805) );
  AND2X1 U1638 ( .A(fifo_array[23]), .B(n4757), .Y(n178) );
  INVX1 U1640 ( .A(n178), .Y(n2806) );
  AND2X1 U1642 ( .A(fifo_array[1079]), .B(n4695), .Y(n1277) );
  INVX1 U1644 ( .A(n1277), .Y(n2807) );
  AND2X1 U1646 ( .A(fifo_array[1046]), .B(n4697), .Y(n1243) );
  INVX1 U1648 ( .A(n1243), .Y(n2808) );
  AND2X1 U1650 ( .A(fifo_array[1006]), .B(n4698), .Y(n1202) );
  INVX1 U1652 ( .A(n1202), .Y(n2809) );
  AND2X1 U1654 ( .A(fifo_array[994]), .B(n4699), .Y(n1190) );
  INVX1 U1656 ( .A(n1190), .Y(n2810) );
  AND2X1 U1658 ( .A(fifo_array[973]), .B(n4700), .Y(n1168) );
  INVX1 U1660 ( .A(n1168), .Y(n2811) );
  AND2X1 U1662 ( .A(fifo_array[962]), .B(n4701), .Y(n1157) );
  INVX1 U1664 ( .A(n1157), .Y(n2812) );
  AND2X1 U1666 ( .A(fifo_array[940]), .B(n4702), .Y(n1134) );
  INVX1 U1668 ( .A(n1134), .Y(n2813) );
  AND2X1 U1670 ( .A(fifo_array[929]), .B(n4703), .Y(n1123) );
  INVX1 U1672 ( .A(n1123), .Y(n2814) );
  AND2X1 U1674 ( .A(fifo_array[913]), .B(n4705), .Y(n1106) );
  INVX1 U1676 ( .A(n1106), .Y(n2815) );
  AND2X1 U1678 ( .A(fifo_array[896]), .B(n4705), .Y(n1089) );
  INVX1 U1680 ( .A(n1089), .Y(n2816) );
  AND2X1 U1682 ( .A(fifo_array[869]), .B(n4707), .Y(n1061) );
  INVX1 U1684 ( .A(n1061), .Y(n2817) );
  AND2X1 U1686 ( .A(fifo_array[857]), .B(n4706), .Y(n1049) );
  INVX1 U1688 ( .A(n1049), .Y(n2818) );
  AND2X1 U1690 ( .A(fifo_array[825]), .B(n4709), .Y(n1015) );
  INVX1 U1691 ( .A(n1015), .Y(n2819) );
  AND2X1 U1693 ( .A(fifo_array[816]), .B(n4708), .Y(n1006) );
  INVX1 U1695 ( .A(n1006), .Y(n2820) );
  AND2X1 U1697 ( .A(fifo_array[795]), .B(n4711), .Y(n984) );
  INVX1 U1699 ( .A(n984), .Y(n2821) );
  AND2X1 U1701 ( .A(fifo_array[783]), .B(n4711), .Y(n972) );
  INVX1 U1703 ( .A(n972), .Y(n2822) );
  AND2X1 U1705 ( .A(fifo_array[762]), .B(n4713), .Y(n950) );
  INVX1 U1707 ( .A(n950), .Y(n2823) );
  AND2X1 U1709 ( .A(fifo_array[750]), .B(n4713), .Y(n938) );
  INVX1 U1711 ( .A(n938), .Y(n2824) );
  AND2X1 U1713 ( .A(fifo_array[729]), .B(n4715), .Y(n916) );
  INVX1 U1715 ( .A(n916), .Y(n2825) );
  AND2X1 U1717 ( .A(fifo_array[717]), .B(n4715), .Y(n904) );
  INVX1 U1719 ( .A(n904), .Y(n2826) );
  AND2X1 U1721 ( .A(fifo_array[703]), .B(n4717), .Y(n889) );
  INVX1 U1723 ( .A(n889), .Y(n2827) );
  AND2X1 U1725 ( .A(fifo_array[670]), .B(n4719), .Y(n855) );
  INVX1 U1727 ( .A(n855), .Y(n2828) );
  AND2X1 U1729 ( .A(fifo_array[637]), .B(n4721), .Y(n821) );
  INVX1 U1731 ( .A(n821), .Y(n2829) );
  AND2X1 U1733 ( .A(fifo_array[604]), .B(n4723), .Y(n787) );
  INVX1 U1735 ( .A(n787), .Y(n2830) );
  AND2X1 U1737 ( .A(fifo_array[564]), .B(n4724), .Y(n745) );
  INVX1 U1739 ( .A(n745), .Y(n2831) );
  AND2X1 U1741 ( .A(fifo_array[552]), .B(n4724), .Y(n733) );
  INVX1 U1743 ( .A(n733), .Y(n2832) );
  AND2X1 U1745 ( .A(fifo_array[531]), .B(n4726), .Y(n711) );
  INVX1 U1747 ( .A(n711), .Y(n2833) );
  AND2X1 U1749 ( .A(fifo_array[520]), .B(n4727), .Y(n700) );
  INVX1 U1751 ( .A(n700), .Y(n2834) );
  AND2X1 U1753 ( .A(fifo_array[498]), .B(n4728), .Y(n677) );
  INVX1 U1755 ( .A(n677), .Y(n2835) );
  AND2X1 U1757 ( .A(fifo_array[487]), .B(n4729), .Y(n666) );
  INVX1 U1759 ( .A(n666), .Y(n2836) );
  AND2X1 U1760 ( .A(fifo_array[471]), .B(n4730), .Y(n649) );
  INVX1 U1763 ( .A(n649), .Y(n2837) );
  AND2X1 U1765 ( .A(fifo_array[454]), .B(n4731), .Y(n632) );
  INVX1 U1767 ( .A(n632), .Y(n2838) );
  AND2X1 U1769 ( .A(fifo_array[427]), .B(n4733), .Y(n604) );
  INVX1 U1771 ( .A(n604), .Y(n2839) );
  AND2X1 U1773 ( .A(fifo_array[415]), .B(n4733), .Y(n592) );
  INVX1 U1775 ( .A(n592), .Y(n2840) );
  AND2X1 U1777 ( .A(fifo_array[383]), .B(n4735), .Y(n559) );
  INVX1 U1779 ( .A(n559), .Y(n2841) );
  AND2X1 U1781 ( .A(fifo_array[374]), .B(n4735), .Y(n550) );
  INVX1 U1783 ( .A(n550), .Y(n2842) );
  AND2X1 U1785 ( .A(fifo_array[353]), .B(n4737), .Y(n528) );
  INVX1 U1787 ( .A(n528), .Y(n2843) );
  AND2X1 U1789 ( .A(fifo_array[341]), .B(n4737), .Y(n516) );
  INVX1 U1791 ( .A(n516), .Y(n2844) );
  AND2X1 U1793 ( .A(fifo_array[320]), .B(n4739), .Y(n494) );
  INVX1 U1795 ( .A(n494), .Y(n2845) );
  AND2X1 U1797 ( .A(fifo_array[308]), .B(n4739), .Y(n482) );
  INVX1 U1799 ( .A(n482), .Y(n2846) );
  AND2X1 U1801 ( .A(fifo_array[287]), .B(n4741), .Y(n459) );
  INVX1 U1803 ( .A(n459), .Y(n2847) );
  AND2X1 U1805 ( .A(fifo_array[275]), .B(n4741), .Y(n447) );
  INVX1 U1807 ( .A(n447), .Y(n2848) );
  AND2X1 U1809 ( .A(fifo_array[261]), .B(n4743), .Y(n431) );
  INVX1 U1811 ( .A(n431), .Y(n2849) );
  AND2X1 U1813 ( .A(fifo_array[228]), .B(n4745), .Y(n396) );
  INVX1 U1815 ( .A(n396), .Y(n2850) );
  AND2X1 U1817 ( .A(fifo_array[195]), .B(n4747), .Y(n361) );
  INVX1 U1819 ( .A(n361), .Y(n2851) );
  AND2X1 U1821 ( .A(fifo_array[162]), .B(n4749), .Y(n326) );
  INVX1 U1823 ( .A(n326), .Y(n2852) );
  AND2X1 U1825 ( .A(fifo_array[122]), .B(n4750), .Y(n284) );
  INVX1 U1827 ( .A(n284), .Y(n2853) );
  AND2X1 U1829 ( .A(fifo_array[110]), .B(n4751), .Y(n272) );
  INVX1 U1830 ( .A(n272), .Y(n2854) );
  AND2X1 U1833 ( .A(fifo_array[89]), .B(n4752), .Y(n249) );
  INVX1 U1835 ( .A(n249), .Y(n2855) );
  AND2X1 U1837 ( .A(fifo_array[78]), .B(n4753), .Y(n238) );
  INVX1 U1839 ( .A(n238), .Y(n2856) );
  AND2X1 U1841 ( .A(fifo_array[56]), .B(n4754), .Y(n214) );
  INVX1 U1843 ( .A(n214), .Y(n2857) );
  AND2X1 U1845 ( .A(fifo_array[45]), .B(n4755), .Y(n203) );
  INVX1 U1847 ( .A(n203), .Y(n2858) );
  AND2X1 U1849 ( .A(fifo_array[29]), .B(n4757), .Y(n184) );
  INVX1 U1851 ( .A(n184), .Y(n2859) );
  AND2X1 U1853 ( .A(fifo_array[12]), .B(n4757), .Y(n167) );
  INVX1 U1855 ( .A(n167), .Y(n2860) );
  AND2X1 U1857 ( .A(fifo_array[1080]), .B(n4695), .Y(n1278) );
  INVX1 U1859 ( .A(n1278), .Y(n2861) );
  AND2X1 U1861 ( .A(fifo_array[1045]), .B(n4697), .Y(n1242) );
  INVX1 U1863 ( .A(n1242), .Y(n2862) );
  AND2X1 U1865 ( .A(fifo_array[1007]), .B(n4698), .Y(n1203) );
  INVX1 U1867 ( .A(n1203), .Y(n2863) );
  AND2X1 U1869 ( .A(fifo_array[996]), .B(n4699), .Y(n1192) );
  INVX1 U1871 ( .A(n1192), .Y(n2864) );
  AND2X1 U1873 ( .A(fifo_array[972]), .B(n4700), .Y(n1167) );
  INVX1 U1875 ( .A(n1167), .Y(n2865) );
  AND2X1 U1877 ( .A(fifo_array[960]), .B(n4701), .Y(n1155) );
  INVX1 U1879 ( .A(n1155), .Y(n2866) );
  AND2X1 U1881 ( .A(fifo_array[947]), .B(n4703), .Y(n1141) );
  INVX1 U1883 ( .A(n1141), .Y(n2867) );
  AND2X1 U1885 ( .A(fifo_array[930]), .B(n4703), .Y(n1124) );
  INVX1 U1887 ( .A(n1124), .Y(n2868) );
  AND2X1 U1889 ( .A(fifo_array[906]), .B(n4704), .Y(n1099) );
  INVX1 U1891 ( .A(n1099), .Y(n2869) );
  AND2X1 U1893 ( .A(fifo_array[895]), .B(n4705), .Y(n1088) );
  INVX1 U1895 ( .A(n1088), .Y(n2870) );
  AND2X1 U1897 ( .A(fifo_array[868]), .B(n4707), .Y(n1060) );
  INVX1 U1899 ( .A(n1060), .Y(n2871) );
  AND2X1 U1900 ( .A(fifo_array[856]), .B(n4706), .Y(n1048) );
  INVX1 U1903 ( .A(n1048), .Y(n2872) );
  AND2X1 U1905 ( .A(fifo_array[829]), .B(n4709), .Y(n1019) );
  INVX1 U1907 ( .A(n1019), .Y(n2873) );
  AND2X1 U1909 ( .A(fifo_array[817]), .B(n4708), .Y(n1007) );
  INVX1 U1911 ( .A(n1007), .Y(n2874) );
  AND2X1 U1913 ( .A(fifo_array[791]), .B(n4711), .Y(n980) );
  INVX1 U1915 ( .A(n980), .Y(n2875) );
  AND2X1 U1917 ( .A(fifo_array[782]), .B(n4711), .Y(n971) );
  INVX1 U1919 ( .A(n971), .Y(n2876) );
  AND2X1 U1921 ( .A(fifo_array[763]), .B(n4713), .Y(n951) );
  INVX1 U1923 ( .A(n951), .Y(n2877) );
  AND2X1 U1925 ( .A(fifo_array[751]), .B(n4713), .Y(n939) );
  INVX1 U1927 ( .A(n939), .Y(n2878) );
  AND2X1 U1929 ( .A(fifo_array[728]), .B(n4715), .Y(n915) );
  INVX1 U1931 ( .A(n915), .Y(n2879) );
  AND2X1 U1933 ( .A(fifo_array[716]), .B(n4715), .Y(n903) );
  INVX1 U1935 ( .A(n903), .Y(n2880) );
  AND2X1 U1937 ( .A(fifo_array[704]), .B(n4717), .Y(n890) );
  INVX1 U1939 ( .A(n890), .Y(n2881) );
  AND2X1 U1941 ( .A(fifo_array[669]), .B(n4719), .Y(n854) );
  INVX1 U1943 ( .A(n854), .Y(n2882) );
  AND2X1 U1945 ( .A(fifo_array[638]), .B(n4721), .Y(n822) );
  INVX1 U1947 ( .A(n822), .Y(n2883) );
  AND2X1 U1949 ( .A(fifo_array[603]), .B(n4723), .Y(n786) );
  INVX1 U1951 ( .A(n786), .Y(n2884) );
  AND2X1 U1953 ( .A(fifo_array[565]), .B(n4724), .Y(n746) );
  INVX1 U1955 ( .A(n746), .Y(n2885) );
  AND2X1 U1957 ( .A(fifo_array[554]), .B(n4725), .Y(n735) );
  INVX1 U1959 ( .A(n735), .Y(n2886) );
  AND2X1 U1961 ( .A(fifo_array[530]), .B(n4726), .Y(n710) );
  INVX1 U1963 ( .A(n710), .Y(n2887) );
  AND2X1 U1965 ( .A(fifo_array[518]), .B(n4726), .Y(n698) );
  INVX1 U1967 ( .A(n698), .Y(n2888) );
  AND2X1 U1969 ( .A(fifo_array[505]), .B(n4728), .Y(n684) );
  INVX1 U1970 ( .A(n684), .Y(n2889) );
  AND2X1 U1973 ( .A(fifo_array[488]), .B(n4729), .Y(n667) );
  INVX1 U1975 ( .A(n667), .Y(n2890) );
  AND2X1 U1977 ( .A(fifo_array[464]), .B(n4730), .Y(n642) );
  INVX1 U1979 ( .A(n642), .Y(n2891) );
  AND2X1 U1981 ( .A(fifo_array[453]), .B(n4731), .Y(n631) );
  INVX1 U1983 ( .A(n631), .Y(n2892) );
  AND2X1 U1985 ( .A(fifo_array[426]), .B(n4733), .Y(n603) );
  INVX1 U1987 ( .A(n603), .Y(n2893) );
  AND2X1 U1989 ( .A(fifo_array[414]), .B(n4733), .Y(n591) );
  INVX1 U1991 ( .A(n591), .Y(n2894) );
  AND2X1 U1993 ( .A(fifo_array[387]), .B(n4735), .Y(n563) );
  INVX1 U1995 ( .A(n563), .Y(n2895) );
  AND2X1 U1997 ( .A(fifo_array[375]), .B(n4735), .Y(n551) );
  INVX1 U1999 ( .A(n551), .Y(n2896) );
  AND2X1 U2001 ( .A(fifo_array[349]), .B(n4737), .Y(n524) );
  INVX1 U2003 ( .A(n524), .Y(n2897) );
  AND2X1 U2005 ( .A(fifo_array[340]), .B(n4737), .Y(n515) );
  INVX1 U2007 ( .A(n515), .Y(n2898) );
  AND2X1 U2009 ( .A(fifo_array[321]), .B(n4739), .Y(n495) );
  INVX1 U2011 ( .A(n495), .Y(n2899) );
  AND2X1 U2013 ( .A(fifo_array[309]), .B(n4739), .Y(n483) );
  INVX1 U2015 ( .A(n483), .Y(n2900) );
  AND2X1 U2017 ( .A(fifo_array[286]), .B(n4741), .Y(n458) );
  INVX1 U2019 ( .A(n458), .Y(n2901) );
  AND2X1 U2021 ( .A(fifo_array[274]), .B(n4741), .Y(n446) );
  INVX1 U2023 ( .A(n446), .Y(n2902) );
  AND2X1 U2025 ( .A(fifo_array[262]), .B(n4743), .Y(n432) );
  INVX1 U2027 ( .A(n432), .Y(n2903) );
  AND2X1 U2029 ( .A(fifo_array[227]), .B(n4745), .Y(n395) );
  INVX1 U2031 ( .A(n395), .Y(n2904) );
  AND2X1 U2033 ( .A(fifo_array[196]), .B(n4747), .Y(n362) );
  INVX1 U2035 ( .A(n362), .Y(n2905) );
  AND2X1 U2037 ( .A(fifo_array[161]), .B(n4749), .Y(n325) );
  INVX1 U2039 ( .A(n325), .Y(n2906) );
  AND2X1 U2040 ( .A(fifo_array[123]), .B(n4751), .Y(n285) );
  INVX1 U2043 ( .A(n285), .Y(n2907) );
  AND2X1 U2045 ( .A(fifo_array[112]), .B(n4751), .Y(n274) );
  INVX1 U2047 ( .A(n274), .Y(n2908) );
  AND2X1 U2049 ( .A(fifo_array[88]), .B(n4753), .Y(n248) );
  INVX1 U2051 ( .A(n248), .Y(n2909) );
  AND2X1 U2053 ( .A(fifo_array[76]), .B(n4753), .Y(n236) );
  INVX1 U2055 ( .A(n236), .Y(n2910) );
  AND2X1 U2057 ( .A(fifo_array[63]), .B(n4755), .Y(n221) );
  INVX1 U2059 ( .A(n221), .Y(n2911) );
  AND2X1 U2061 ( .A(fifo_array[46]), .B(n4755), .Y(n204) );
  INVX1 U2063 ( .A(n204), .Y(n2912) );
  AND2X1 U2065 ( .A(fifo_array[22]), .B(n4756), .Y(n177) );
  INVX1 U2067 ( .A(n177), .Y(n2913) );
  AND2X1 U2069 ( .A(fifo_array[11]), .B(n4757), .Y(n166) );
  INVX1 U2071 ( .A(n166), .Y(n2914) );
  AND2X1 U2073 ( .A(fifo_array[1077]), .B(n4695), .Y(n1275) );
  INVX1 U2075 ( .A(n1275), .Y(n2915) );
  AND2X1 U2077 ( .A(fifo_array[1044]), .B(n4697), .Y(n1241) );
  INVX1 U2079 ( .A(n1241), .Y(n2916) );
  AND2X1 U2081 ( .A(fifo_array[1008]), .B(n4698), .Y(n1204) );
  INVX1 U2083 ( .A(n1204), .Y(n2917) );
  AND2X1 U2085 ( .A(fifo_array[997]), .B(n4699), .Y(n1193) );
  INVX1 U2087 ( .A(n1193), .Y(n2918) );
  AND2X1 U2089 ( .A(fifo_array[981]), .B(n4701), .Y(n1176) );
  INVX1 U2091 ( .A(n1176), .Y(n2919) );
  AND2X1 U2093 ( .A(fifo_array[964]), .B(n4701), .Y(n1159) );
  INVX1 U2095 ( .A(n1159), .Y(n2920) );
  AND2X1 U2097 ( .A(fifo_array[938]), .B(n4702), .Y(n1132) );
  INVX1 U2099 ( .A(n1132), .Y(n2921) );
  AND2X1 U2101 ( .A(fifo_array[926]), .B(n4703), .Y(n1120) );
  INVX1 U2103 ( .A(n1120), .Y(n2922) );
  AND2X1 U2105 ( .A(fifo_array[905]), .B(n4704), .Y(n1098) );
  INVX1 U2107 ( .A(n1098), .Y(n2923) );
  AND2X1 U2109 ( .A(fifo_array[894]), .B(n4705), .Y(n1087) );
  INVX1 U2110 ( .A(n1087), .Y(n2924) );
  AND2X1 U2113 ( .A(fifo_array[867]), .B(n4707), .Y(n1059) );
  INVX1 U2115 ( .A(n1059), .Y(n2925) );
  AND2X1 U2117 ( .A(fifo_array[855]), .B(n4707), .Y(n1047) );
  INVX1 U2119 ( .A(n1047), .Y(n2926) );
  AND2X1 U2121 ( .A(fifo_array[830]), .B(n4709), .Y(n1020) );
  INVX1 U2123 ( .A(n1020), .Y(n2927) );
  AND2X1 U2125 ( .A(fifo_array[818]), .B(n4709), .Y(n1008) );
  INVX1 U2127 ( .A(n1008), .Y(n2928) );
  AND2X1 U2129 ( .A(fifo_array[797]), .B(n4711), .Y(n986) );
  INVX1 U2131 ( .A(n986), .Y(n2929) );
  AND2X1 U2133 ( .A(fifo_array[785]), .B(n4711), .Y(n974) );
  INVX1 U2135 ( .A(n974), .Y(n2930) );
  AND2X1 U2137 ( .A(fifo_array[757]), .B(n4713), .Y(n945) );
  INVX1 U2139 ( .A(n945), .Y(n2931) );
  AND2X1 U2141 ( .A(fifo_array[748]), .B(n4713), .Y(n936) );
  INVX1 U2143 ( .A(n936), .Y(n2932) );
  AND2X1 U2145 ( .A(fifo_array[727]), .B(n4715), .Y(n914) );
  INVX1 U2147 ( .A(n914), .Y(n2933) );
  AND2X1 U2149 ( .A(fifo_array[715]), .B(n4715), .Y(n902) );
  INVX1 U2151 ( .A(n902), .Y(n2934) );
  AND2X1 U2153 ( .A(fifo_array[705]), .B(n4717), .Y(n891) );
  INVX1 U2155 ( .A(n891), .Y(n2935) );
  AND2X1 U2157 ( .A(fifo_array[672]), .B(n4719), .Y(n857) );
  INVX1 U2159 ( .A(n857), .Y(n2936) );
  AND2X1 U2161 ( .A(fifo_array[635]), .B(n4721), .Y(n819) );
  INVX1 U2163 ( .A(n819), .Y(n2937) );
  AND2X1 U2165 ( .A(fifo_array[602]), .B(n4723), .Y(n785) );
  INVX1 U2167 ( .A(n785), .Y(n2938) );
  AND2X1 U2169 ( .A(fifo_array[566]), .B(n4724), .Y(n747) );
  INVX1 U2171 ( .A(n747), .Y(n2939) );
  AND2X1 U2173 ( .A(fifo_array[555]), .B(n4725), .Y(n736) );
  INVX1 U2175 ( .A(n736), .Y(n2940) );
  AND2X1 U2177 ( .A(fifo_array[539]), .B(n4727), .Y(n719) );
  INVX1 U2179 ( .A(n719), .Y(n2941) );
  AND2X1 U2180 ( .A(fifo_array[522]), .B(n4727), .Y(n702) );
  INVX1 U2183 ( .A(n702), .Y(n2942) );
  AND2X1 U2185 ( .A(fifo_array[496]), .B(n4728), .Y(n675) );
  INVX1 U2187 ( .A(n675), .Y(n2943) );
  AND2X1 U2189 ( .A(fifo_array[484]), .B(n4729), .Y(n663) );
  INVX1 U2191 ( .A(n663), .Y(n2944) );
  AND2X1 U2193 ( .A(fifo_array[463]), .B(n4730), .Y(n641) );
  INVX1 U2195 ( .A(n641), .Y(n2945) );
  AND2X1 U2197 ( .A(fifo_array[452]), .B(n4731), .Y(n630) );
  INVX1 U2199 ( .A(n630), .Y(n2946) );
  AND2X1 U2201 ( .A(fifo_array[425]), .B(n4733), .Y(n602) );
  INVX1 U2203 ( .A(n602), .Y(n2947) );
  AND2X1 U2205 ( .A(fifo_array[413]), .B(n4733), .Y(n590) );
  INVX1 U2207 ( .A(n590), .Y(n2948) );
  AND2X1 U2209 ( .A(fifo_array[388]), .B(n4735), .Y(n564) );
  INVX1 U2211 ( .A(n564), .Y(n2949) );
  AND2X1 U2213 ( .A(fifo_array[376]), .B(n4735), .Y(n552) );
  INVX1 U2215 ( .A(n552), .Y(n2950) );
  AND2X1 U2217 ( .A(fifo_array[355]), .B(n4737), .Y(n530) );
  INVX1 U2219 ( .A(n530), .Y(n2951) );
  AND2X1 U2221 ( .A(fifo_array[343]), .B(n4737), .Y(n518) );
  INVX1 U2223 ( .A(n518), .Y(n2952) );
  AND2X1 U2225 ( .A(fifo_array[315]), .B(n4739), .Y(n489) );
  INVX1 U2227 ( .A(n489), .Y(n2953) );
  AND2X1 U2229 ( .A(fifo_array[306]), .B(n4739), .Y(n480) );
  INVX1 U2231 ( .A(n480), .Y(n2954) );
  AND2X1 U2233 ( .A(fifo_array[285]), .B(n4741), .Y(n457) );
  INVX1 U2235 ( .A(n457), .Y(n2955) );
  AND2X1 U2237 ( .A(fifo_array[273]), .B(n4741), .Y(n445) );
  INVX1 U2239 ( .A(n445), .Y(n2956) );
  AND2X1 U2241 ( .A(fifo_array[263]), .B(n4743), .Y(n433) );
  INVX1 U2243 ( .A(n433), .Y(n2957) );
  AND2X1 U2245 ( .A(fifo_array[230]), .B(n4745), .Y(n398) );
  INVX1 U2247 ( .A(n398), .Y(n2958) );
  AND2X1 U2249 ( .A(fifo_array[193]), .B(n4747), .Y(n359) );
  INVX1 U2250 ( .A(n359), .Y(n2959) );
  AND2X1 U2253 ( .A(fifo_array[160]), .B(n4749), .Y(n324) );
  INVX1 U2255 ( .A(n324), .Y(n2960) );
  AND2X1 U2257 ( .A(fifo_array[124]), .B(n4751), .Y(n286) );
  INVX1 U2259 ( .A(n286), .Y(n2961) );
  AND2X1 U2261 ( .A(fifo_array[113]), .B(n4751), .Y(n275) );
  INVX1 U2263 ( .A(n275), .Y(n2962) );
  AND2X1 U2265 ( .A(fifo_array[97]), .B(n4753), .Y(n257) );
  INVX1 U2267 ( .A(n257), .Y(n2963) );
  AND2X1 U2269 ( .A(fifo_array[80]), .B(n4753), .Y(n240) );
  INVX1 U2271 ( .A(n240), .Y(n2964) );
  AND2X1 U2273 ( .A(fifo_array[54]), .B(n4755), .Y(n212) );
  INVX1 U2275 ( .A(n212), .Y(n2965) );
  AND2X1 U2277 ( .A(fifo_array[42]), .B(n4755), .Y(n200) );
  INVX1 U2279 ( .A(n200), .Y(n2966) );
  AND2X1 U2281 ( .A(fifo_array[21]), .B(n4756), .Y(n176) );
  INVX1 U2283 ( .A(n176), .Y(n2967) );
  AND2X1 U2285 ( .A(fifo_array[10]), .B(n4757), .Y(n165) );
  INVX1 U2287 ( .A(n165), .Y(n2968) );
  AND2X1 U2289 ( .A(fifo_array[1078]), .B(n4695), .Y(n1276) );
  INVX1 U2291 ( .A(n1276), .Y(n2969) );
  AND2X1 U2293 ( .A(fifo_array[1043]), .B(n4697), .Y(n1240) );
  INVX1 U2295 ( .A(n1240), .Y(n2970) );
  AND2X1 U2297 ( .A(fifo_array[1015]), .B(n4699), .Y(n1211) );
  INVX1 U2299 ( .A(n1211), .Y(n2971) );
  AND2X1 U2301 ( .A(fifo_array[998]), .B(n4699), .Y(n1194) );
  INVX1 U2303 ( .A(n1194), .Y(n2972) );
  AND2X1 U2305 ( .A(fifo_array[974]), .B(n4700), .Y(n1169) );
  INVX1 U2307 ( .A(n1169), .Y(n2973) );
  AND2X1 U2309 ( .A(fifo_array[963]), .B(n4701), .Y(n1158) );
  INVX1 U2311 ( .A(n1158), .Y(n2974) );
  AND2X1 U2313 ( .A(fifo_array[939]), .B(n4702), .Y(n1133) );
  INVX1 U2315 ( .A(n1133), .Y(n2975) );
  AND2X1 U2317 ( .A(fifo_array[928]), .B(n4703), .Y(n1122) );
  INVX1 U2319 ( .A(n1122), .Y(n2976) );
  AND2X1 U2320 ( .A(fifo_array[904]), .B(n4704), .Y(n1097) );
  INVX1 U2324 ( .A(n1097), .Y(n2977) );
  AND2X1 U2326 ( .A(fifo_array[892]), .B(n4705), .Y(n1085) );
  INVX1 U2328 ( .A(n1085), .Y(n2978) );
  AND2X1 U2330 ( .A(fifo_array[866]), .B(n4707), .Y(n1058) );
  INVX1 U2332 ( .A(n1058), .Y(n2979) );
  AND2X1 U2333 ( .A(fifo_array[854]), .B(n4706), .Y(n1046) );
  INVX1 U2334 ( .A(n1046), .Y(n2980) );
  AND2X1 U2384 ( .A(fifo_array[831]), .B(n4709), .Y(n1021) );
  INVX1 U2386 ( .A(n1021), .Y(n2981) );
  AND2X1 U2390 ( .A(fifo_array[819]), .B(n4708), .Y(n1009) );
  INVX1 U2393 ( .A(n1009), .Y(n2982) );
  AND2X1 U2395 ( .A(fifo_array[796]), .B(n4711), .Y(n985) );
  INVX1 U2400 ( .A(n985), .Y(n2983) );
  AND2X1 U2401 ( .A(fifo_array[784]), .B(n4711), .Y(n973) );
  INVX1 U2403 ( .A(n973), .Y(n2984) );
  AND2X1 U2404 ( .A(fifo_array[761]), .B(n4713), .Y(n949) );
  INVX1 U2405 ( .A(n949), .Y(n2985) );
  AND2X1 U2406 ( .A(fifo_array[749]), .B(n4713), .Y(n937) );
  INVX1 U2407 ( .A(n937), .Y(n2986) );
  AND2X1 U2408 ( .A(fifo_array[723]), .B(n4715), .Y(n910) );
  INVX1 U2409 ( .A(n910), .Y(n2987) );
  AND2X1 U2410 ( .A(fifo_array[714]), .B(n4715), .Y(n901) );
  INVX1 U2411 ( .A(n901), .Y(n2988) );
  AND2X1 U2412 ( .A(fifo_array[706]), .B(n4717), .Y(n892) );
  INVX1 U2413 ( .A(n892), .Y(n2989) );
  AND2X1 U2414 ( .A(fifo_array[671]), .B(n4719), .Y(n856) );
  INVX1 U2415 ( .A(n856), .Y(n2990) );
  AND2X1 U2416 ( .A(fifo_array[636]), .B(n4721), .Y(n820) );
  INVX1 U2417 ( .A(n820), .Y(n2991) );
  AND2X1 U2418 ( .A(fifo_array[601]), .B(n4723), .Y(n784) );
  INVX1 U2419 ( .A(n784), .Y(n2992) );
  AND2X1 U2420 ( .A(fifo_array[573]), .B(n4725), .Y(n754) );
  INVX1 U2421 ( .A(n754), .Y(n2993) );
  AND2X1 U2422 ( .A(fifo_array[556]), .B(n4725), .Y(n737) );
  INVX1 U2423 ( .A(n737), .Y(n2994) );
  AND2X1 U2424 ( .A(fifo_array[532]), .B(n4726), .Y(n712) );
  INVX1 U2425 ( .A(n712), .Y(n2995) );
  AND2X1 U2426 ( .A(fifo_array[521]), .B(n4727), .Y(n701) );
  INVX1 U2427 ( .A(n701), .Y(n2996) );
  AND2X1 U2428 ( .A(fifo_array[497]), .B(n4728), .Y(n676) );
  INVX1 U2429 ( .A(n676), .Y(n2997) );
  AND2X1 U2430 ( .A(fifo_array[486]), .B(n4729), .Y(n665) );
  INVX1 U2431 ( .A(n665), .Y(n2998) );
  AND2X1 U2432 ( .A(fifo_array[462]), .B(n4730), .Y(n640) );
  INVX1 U2433 ( .A(n640), .Y(n2999) );
  AND2X1 U2434 ( .A(fifo_array[450]), .B(n4731), .Y(n628) );
  INVX1 U2435 ( .A(n628), .Y(n3000) );
  AND2X1 U2436 ( .A(fifo_array[424]), .B(n4733), .Y(n601) );
  INVX1 U2437 ( .A(n601), .Y(n3001) );
  AND2X1 U2438 ( .A(fifo_array[412]), .B(n4733), .Y(n589) );
  INVX1 U2439 ( .A(n589), .Y(n3002) );
  AND2X1 U2440 ( .A(fifo_array[389]), .B(n4735), .Y(n565) );
  INVX1 U2441 ( .A(n565), .Y(n3003) );
  AND2X1 U2442 ( .A(fifo_array[377]), .B(n4735), .Y(n553) );
  INVX1 U2443 ( .A(n553), .Y(n3004) );
  AND2X1 U2444 ( .A(fifo_array[354]), .B(n4737), .Y(n529) );
  INVX1 U2445 ( .A(n529), .Y(n3005) );
  AND2X1 U2446 ( .A(fifo_array[342]), .B(n4737), .Y(n517) );
  INVX1 U2447 ( .A(n517), .Y(n3006) );
  AND2X1 U2448 ( .A(fifo_array[319]), .B(n4739), .Y(n493) );
  INVX1 U2449 ( .A(n493), .Y(n3007) );
  AND2X1 U2450 ( .A(fifo_array[307]), .B(n4739), .Y(n481) );
  INVX1 U2451 ( .A(n481), .Y(n3008) );
  AND2X1 U2452 ( .A(fifo_array[281]), .B(n4741), .Y(n453) );
  INVX1 U2453 ( .A(n453), .Y(n3009) );
  AND2X1 U2454 ( .A(fifo_array[272]), .B(n4741), .Y(n444) );
  INVX1 U2455 ( .A(n444), .Y(n3010) );
  AND2X1 U2456 ( .A(fifo_array[264]), .B(n4743), .Y(n434) );
  INVX1 U2457 ( .A(n434), .Y(n3011) );
  AND2X1 U2458 ( .A(fifo_array[229]), .B(n4745), .Y(n397) );
  INVX1 U2459 ( .A(n397), .Y(n3012) );
  AND2X1 U2460 ( .A(fifo_array[194]), .B(n4747), .Y(n360) );
  INVX1 U2461 ( .A(n360), .Y(n3013) );
  AND2X1 U2462 ( .A(fifo_array[159]), .B(n4749), .Y(n323) );
  INVX1 U2463 ( .A(n323), .Y(n3014) );
  AND2X1 U2464 ( .A(fifo_array[131]), .B(n4751), .Y(n293) );
  INVX1 U2465 ( .A(n293), .Y(n3015) );
  AND2X1 U2466 ( .A(fifo_array[114]), .B(n4751), .Y(n276) );
  INVX1 U2467 ( .A(n276), .Y(n3016) );
  AND2X1 U2468 ( .A(fifo_array[90]), .B(n4753), .Y(n250) );
  INVX1 U2469 ( .A(n250), .Y(n3017) );
  AND2X1 U2470 ( .A(fifo_array[79]), .B(n4753), .Y(n239) );
  INVX1 U2471 ( .A(n239), .Y(n3018) );
  AND2X1 U2472 ( .A(fifo_array[55]), .B(n4755), .Y(n213) );
  INVX1 U2473 ( .A(n213), .Y(n3019) );
  AND2X1 U2474 ( .A(fifo_array[44]), .B(n4755), .Y(n202) );
  INVX1 U2475 ( .A(n202), .Y(n3020) );
  AND2X1 U2476 ( .A(fifo_array[20]), .B(n4757), .Y(n175) );
  INVX1 U2477 ( .A(n175), .Y(n3021) );
  AND2X1 U2478 ( .A(fifo_array[8]), .B(n4757), .Y(n163) );
  INVX1 U2479 ( .A(n163), .Y(n3022) );
  AND2X1 U2480 ( .A(n4808), .B(n3457), .Y(n1292) );
  INVX1 U2481 ( .A(n1292), .Y(n3023) );
  BUFX2 U2482 ( .A(n1302), .Y(n3024) );
  AND2X1 U2483 ( .A(fifo_array[1068]), .B(n4695), .Y(n1266) );
  INVX1 U2484 ( .A(n1266), .Y(n3025) );
  AND2X1 U2485 ( .A(fifo_array[1056]), .B(n4695), .Y(n1254) );
  INVX1 U2486 ( .A(n1254), .Y(n3026) );
  AND2X1 U2487 ( .A(fifo_array[1035]), .B(n4697), .Y(n1232) );
  INVX1 U2488 ( .A(n1232), .Y(n3027) );
  AND2X1 U2489 ( .A(fifo_array[1023]), .B(n4697), .Y(n1220) );
  INVX1 U2490 ( .A(n1220), .Y(n3028) );
  AND2X1 U2491 ( .A(fifo_array[1002]), .B(n4699), .Y(n1198) );
  INVX1 U2492 ( .A(n1198), .Y(n3029) );
  AND2X1 U2493 ( .A(fifo_array[990]), .B(n4699), .Y(n1186) );
  INVX1 U2494 ( .A(n1186), .Y(n3030) );
  AND2X1 U2495 ( .A(fifo_array[969]), .B(n4701), .Y(n1164) );
  INVX1 U2496 ( .A(n1164), .Y(n3031) );
  AND2X1 U2497 ( .A(fifo_array[957]), .B(n4701), .Y(n1152) );
  INVX1 U2498 ( .A(n1152), .Y(n3032) );
  AND2X1 U2499 ( .A(fifo_array[936]), .B(n4703), .Y(n1130) );
  INVX1 U2500 ( .A(n1130), .Y(n3033) );
  AND2X1 U2501 ( .A(fifo_array[924]), .B(n4703), .Y(n1118) );
  INVX1 U2502 ( .A(n1118), .Y(n3034) );
  AND2X1 U2503 ( .A(fifo_array[903]), .B(n4705), .Y(n1096) );
  INVX1 U2504 ( .A(n1096), .Y(n3035) );
  AND2X1 U2505 ( .A(fifo_array[891]), .B(n4705), .Y(n1084) );
  INVX1 U2506 ( .A(n1084), .Y(n3036) );
  AND2X1 U2507 ( .A(fifo_array[879]), .B(n4707), .Y(n1071) );
  INVX1 U2508 ( .A(n1071), .Y(n3037) );
  AND2X1 U2509 ( .A(fifo_array[862]), .B(n4707), .Y(n1054) );
  INVX1 U2510 ( .A(n1054), .Y(n3038) );
  AND2X1 U2511 ( .A(fifo_array[839]), .B(n4709), .Y(n1029) );
  INVX1 U2512 ( .A(n1029), .Y(n3039) );
  AND2X1 U2513 ( .A(fifo_array[806]), .B(n4711), .Y(n995) );
  INVX1 U2514 ( .A(n995), .Y(n3040) );
  AND2X1 U2515 ( .A(fifo_array[773]), .B(n4713), .Y(n961) );
  INVX1 U2516 ( .A(n961), .Y(n3041) );
  AND2X1 U2517 ( .A(fifo_array[740]), .B(n4715), .Y(n927) );
  INVX1 U2518 ( .A(n927), .Y(n3042) );
  AND2X1 U2519 ( .A(fifo_array[689]), .B(n4717), .Y(n875) );
  INVX1 U2520 ( .A(n875), .Y(n3043) );
  AND2X1 U2521 ( .A(fifo_array[680]), .B(n4717), .Y(n866) );
  INVX1 U2522 ( .A(n866), .Y(n3044) );
  AND2X1 U2523 ( .A(fifo_array[659]), .B(n4719), .Y(n844) );
  INVX1 U2524 ( .A(n844), .Y(n3045) );
  AND2X1 U2525 ( .A(fifo_array[647]), .B(n4719), .Y(n832) );
  INVX1 U2526 ( .A(n832), .Y(n3046) );
  AND2X1 U2527 ( .A(fifo_array[626]), .B(n4721), .Y(n810) );
  INVX1 U2528 ( .A(n810), .Y(n3047) );
  AND2X1 U2529 ( .A(fifo_array[614]), .B(n4721), .Y(n798) );
  INVX1 U2530 ( .A(n798), .Y(n3048) );
  AND2X1 U2531 ( .A(fifo_array[593]), .B(n4723), .Y(n776) );
  INVX1 U2532 ( .A(n776), .Y(n3049) );
  AND2X1 U2533 ( .A(fifo_array[581]), .B(n4723), .Y(n764) );
  INVX1 U2534 ( .A(n764), .Y(n3050) );
  AND2X1 U2535 ( .A(fifo_array[560]), .B(n4725), .Y(n741) );
  INVX1 U2536 ( .A(n741), .Y(n3051) );
  AND2X1 U2537 ( .A(fifo_array[548]), .B(n4725), .Y(n729) );
  INVX1 U2538 ( .A(n729), .Y(n3052) );
  AND2X1 U2539 ( .A(fifo_array[527]), .B(n4727), .Y(n707) );
  INVX1 U2540 ( .A(n707), .Y(n3053) );
  AND2X1 U2541 ( .A(fifo_array[515]), .B(n4727), .Y(n695) );
  INVX1 U2542 ( .A(n695), .Y(n3054) );
  AND2X1 U2543 ( .A(fifo_array[494]), .B(n4729), .Y(n673) );
  INVX1 U2544 ( .A(n673), .Y(n3055) );
  AND2X1 U2545 ( .A(fifo_array[482]), .B(n4729), .Y(n661) );
  INVX1 U2546 ( .A(n661), .Y(n3056) );
  AND2X1 U2547 ( .A(fifo_array[461]), .B(n4731), .Y(n639) );
  INVX1 U2548 ( .A(n639), .Y(n3057) );
  AND2X1 U2549 ( .A(fifo_array[449]), .B(n4731), .Y(n627) );
  INVX1 U2550 ( .A(n627), .Y(n3058) );
  AND2X1 U2551 ( .A(fifo_array[437]), .B(n4732), .Y(n614) );
  INVX1 U2552 ( .A(n614), .Y(n3059) );
  AND2X1 U2553 ( .A(fifo_array[420]), .B(n4733), .Y(n597) );
  INVX1 U2554 ( .A(n597), .Y(n3060) );
  AND2X1 U2555 ( .A(fifo_array[397]), .B(n4735), .Y(n573) );
  INVX1 U2556 ( .A(n573), .Y(n3061) );
  AND2X1 U2557 ( .A(fifo_array[364]), .B(n4737), .Y(n539) );
  INVX1 U2558 ( .A(n539), .Y(n3062) );
  AND2X1 U2559 ( .A(fifo_array[331]), .B(n4739), .Y(n505) );
  INVX1 U2560 ( .A(n505), .Y(n3063) );
  AND2X1 U2561 ( .A(fifo_array[298]), .B(n4741), .Y(n470) );
  INVX1 U2562 ( .A(n470), .Y(n3064) );
  AND2X1 U2563 ( .A(fifo_array[247]), .B(n4743), .Y(n417) );
  INVX1 U2564 ( .A(n417), .Y(n3065) );
  AND2X1 U2565 ( .A(fifo_array[238]), .B(n4742), .Y(n408) );
  INVX1 U2566 ( .A(n408), .Y(n3066) );
  AND2X1 U2567 ( .A(fifo_array[217]), .B(n4745), .Y(n385) );
  INVX1 U2568 ( .A(n385), .Y(n3067) );
  AND2X1 U2569 ( .A(fifo_array[205]), .B(n4744), .Y(n373) );
  INVX1 U2570 ( .A(n373), .Y(n3068) );
  AND2X1 U2571 ( .A(fifo_array[184]), .B(n4747), .Y(n350) );
  INVX1 U2572 ( .A(n350), .Y(n3069) );
  AND2X1 U2573 ( .A(fifo_array[172]), .B(n4746), .Y(n338) );
  INVX1 U2574 ( .A(n338), .Y(n3070) );
  AND2X1 U2575 ( .A(fifo_array[151]), .B(n4749), .Y(n315) );
  INVX1 U2576 ( .A(n315), .Y(n3071) );
  AND2X1 U2577 ( .A(fifo_array[139]), .B(n4748), .Y(n303) );
  INVX1 U2578 ( .A(n303), .Y(n3072) );
  AND2X1 U2579 ( .A(fifo_array[118]), .B(n4751), .Y(n280) );
  INVX1 U2580 ( .A(n280), .Y(n3073) );
  AND2X1 U2581 ( .A(fifo_array[106]), .B(n4750), .Y(n268) );
  INVX1 U2582 ( .A(n268), .Y(n3074) );
  AND2X1 U2583 ( .A(fifo_array[85]), .B(n4753), .Y(n245) );
  INVX1 U2584 ( .A(n245), .Y(n3075) );
  AND2X1 U2585 ( .A(fifo_array[73]), .B(n4752), .Y(n233) );
  INVX1 U2586 ( .A(n233), .Y(n3076) );
  AND2X1 U2587 ( .A(fifo_array[52]), .B(n4755), .Y(n210) );
  INVX1 U2588 ( .A(n210), .Y(n3077) );
  AND2X1 U2589 ( .A(fifo_array[40]), .B(n4754), .Y(n198) );
  INVX1 U2590 ( .A(n198), .Y(n3078) );
  AND2X1 U2591 ( .A(fifo_array[19]), .B(n4757), .Y(n174) );
  INVX1 U2592 ( .A(n174), .Y(n3079) );
  AND2X1 U2593 ( .A(fifo_array[7]), .B(n4756), .Y(n162) );
  INVX1 U2594 ( .A(n162), .Y(n3080) );
  AND2X1 U2595 ( .A(n68), .B(n3457), .Y(n1291) );
  INVX1 U2596 ( .A(n1291), .Y(n3081) );
  BUFX2 U2597 ( .A(n1296), .Y(n3082) );
  AND2X1 U2598 ( .A(fifo_array[1069]), .B(n4695), .Y(n1267) );
  INVX1 U2599 ( .A(n1267), .Y(n3083) );
  AND2X1 U2600 ( .A(fifo_array[1057]), .B(n4694), .Y(n1255) );
  INVX1 U2601 ( .A(n1255), .Y(n3084) );
  AND2X1 U2602 ( .A(fifo_array[1034]), .B(n4697), .Y(n1231) );
  INVX1 U2603 ( .A(n1231), .Y(n3085) );
  AND2X1 U2604 ( .A(fifo_array[1022]), .B(n4696), .Y(n1219) );
  INVX1 U2605 ( .A(n1219), .Y(n3086) );
  AND2X1 U2606 ( .A(fifo_array[1003]), .B(n4699), .Y(n1199) );
  INVX1 U2607 ( .A(n1199), .Y(n3087) );
  AND2X1 U2608 ( .A(fifo_array[991]), .B(n4698), .Y(n1187) );
  INVX1 U2609 ( .A(n1187), .Y(n3088) );
  AND2X1 U2610 ( .A(fifo_array[968]), .B(n4701), .Y(n1163) );
  INVX1 U2611 ( .A(n1163), .Y(n3089) );
  AND2X1 U2612 ( .A(fifo_array[956]), .B(n4700), .Y(n1151) );
  INVX1 U2613 ( .A(n1151), .Y(n3090) );
  AND2X1 U2614 ( .A(fifo_array[937]), .B(n4703), .Y(n1131) );
  INVX1 U2615 ( .A(n1131), .Y(n3091) );
  AND2X1 U2616 ( .A(fifo_array[925]), .B(n4702), .Y(n1119) );
  INVX1 U2617 ( .A(n1119), .Y(n3092) );
  AND2X1 U2618 ( .A(fifo_array[902]), .B(n4705), .Y(n1095) );
  INVX1 U2619 ( .A(n1095), .Y(n3093) );
  AND2X1 U2620 ( .A(fifo_array[890]), .B(n4704), .Y(n1083) );
  INVX1 U2621 ( .A(n1083), .Y(n3094) );
  AND2X1 U2622 ( .A(fifo_array[872]), .B(n4706), .Y(n1064) );
  INVX1 U2623 ( .A(n1064), .Y(n3095) );
  AND2X1 U2624 ( .A(fifo_array[861]), .B(n4707), .Y(n1053) );
  INVX1 U2625 ( .A(n1053), .Y(n3096) );
  AND2X1 U2626 ( .A(fifo_array[840]), .B(n4709), .Y(n1030) );
  INVX1 U2627 ( .A(n1030), .Y(n3097) );
  AND2X1 U2628 ( .A(fifo_array[805]), .B(n4711), .Y(n994) );
  INVX1 U2629 ( .A(n994), .Y(n3098) );
  AND2X1 U2630 ( .A(fifo_array[774]), .B(n4713), .Y(n962) );
  INVX1 U2631 ( .A(n962), .Y(n3099) );
  AND2X1 U2632 ( .A(fifo_array[739]), .B(n4715), .Y(n926) );
  INVX1 U2633 ( .A(n926), .Y(n3100) );
  AND2X1 U2634 ( .A(fifo_array[693]), .B(n4717), .Y(n879) );
  INVX1 U2635 ( .A(n879), .Y(n3101) );
  AND2X1 U2636 ( .A(fifo_array[681]), .B(n4716), .Y(n867) );
  INVX1 U2637 ( .A(n867), .Y(n3102) );
  AND2X1 U2638 ( .A(fifo_array[655]), .B(n4719), .Y(n840) );
  INVX1 U2639 ( .A(n840), .Y(n3103) );
  AND2X1 U2640 ( .A(fifo_array[646]), .B(n4718), .Y(n831) );
  INVX1 U2641 ( .A(n831), .Y(n3104) );
  AND2X1 U2642 ( .A(fifo_array[627]), .B(n4721), .Y(n811) );
  INVX1 U2643 ( .A(n811), .Y(n3105) );
  AND2X1 U2644 ( .A(fifo_array[615]), .B(n4720), .Y(n799) );
  INVX1 U2645 ( .A(n799), .Y(n3106) );
  AND2X1 U2646 ( .A(fifo_array[592]), .B(n4723), .Y(n775) );
  INVX1 U2647 ( .A(n775), .Y(n3107) );
  AND2X1 U2648 ( .A(fifo_array[580]), .B(n4722), .Y(n763) );
  INVX1 U2649 ( .A(n763), .Y(n3108) );
  AND2X1 U2650 ( .A(fifo_array[561]), .B(n4725), .Y(n742) );
  INVX1 U2651 ( .A(n742), .Y(n3109) );
  AND2X1 U2652 ( .A(fifo_array[549]), .B(n4724), .Y(n730) );
  INVX1 U2653 ( .A(n730), .Y(n3110) );
  AND2X1 U2654 ( .A(fifo_array[526]), .B(n4727), .Y(n706) );
  INVX1 U2655 ( .A(n706), .Y(n3111) );
  AND2X1 U2656 ( .A(fifo_array[514]), .B(n4726), .Y(n694) );
  INVX1 U2657 ( .A(n694), .Y(n3112) );
  AND2X1 U2658 ( .A(fifo_array[495]), .B(n4729), .Y(n674) );
  INVX1 U2659 ( .A(n674), .Y(n3113) );
  AND2X1 U2660 ( .A(fifo_array[483]), .B(n4728), .Y(n662) );
  INVX1 U2661 ( .A(n662), .Y(n3114) );
  AND2X1 U2662 ( .A(fifo_array[460]), .B(n4731), .Y(n638) );
  INVX1 U2663 ( .A(n638), .Y(n3115) );
  AND2X1 U2664 ( .A(fifo_array[448]), .B(n4730), .Y(n626) );
  INVX1 U2665 ( .A(n626), .Y(n3116) );
  AND2X1 U2666 ( .A(fifo_array[430]), .B(n4732), .Y(n607) );
  INVX1 U2667 ( .A(n607), .Y(n3117) );
  AND2X1 U2668 ( .A(fifo_array[419]), .B(n4733), .Y(n596) );
  INVX1 U2669 ( .A(n596), .Y(n3118) );
  AND2X1 U2670 ( .A(fifo_array[398]), .B(n4735), .Y(n574) );
  INVX1 U2671 ( .A(n574), .Y(n3119) );
  AND2X1 U2672 ( .A(fifo_array[363]), .B(n4737), .Y(n538) );
  INVX1 U2673 ( .A(n538), .Y(n3120) );
  AND2X1 U2674 ( .A(fifo_array[332]), .B(n4739), .Y(n506) );
  INVX1 U2675 ( .A(n506), .Y(n3121) );
  AND2X1 U2676 ( .A(fifo_array[297]), .B(n4741), .Y(n469) );
  INVX1 U2677 ( .A(n469), .Y(n3122) );
  AND2X1 U2678 ( .A(fifo_array[251]), .B(n4743), .Y(n421) );
  INVX1 U2679 ( .A(n421), .Y(n3123) );
  AND2X1 U2680 ( .A(fifo_array[239]), .B(n4743), .Y(n409) );
  INVX1 U2681 ( .A(n409), .Y(n3124) );
  AND2X1 U2682 ( .A(fifo_array[213]), .B(n4745), .Y(n381) );
  INVX1 U2683 ( .A(n381), .Y(n3125) );
  AND2X1 U2684 ( .A(fifo_array[204]), .B(n4745), .Y(n372) );
  INVX1 U2685 ( .A(n372), .Y(n3126) );
  AND2X1 U2686 ( .A(fifo_array[185]), .B(n4747), .Y(n351) );
  INVX1 U2687 ( .A(n351), .Y(n3127) );
  AND2X1 U2688 ( .A(fifo_array[173]), .B(n4747), .Y(n339) );
  INVX1 U2689 ( .A(n339), .Y(n3128) );
  AND2X1 U2690 ( .A(fifo_array[150]), .B(n4749), .Y(n314) );
  INVX1 U2691 ( .A(n314), .Y(n3129) );
  AND2X1 U2692 ( .A(fifo_array[138]), .B(n4749), .Y(n302) );
  INVX1 U2693 ( .A(n302), .Y(n3130) );
  AND2X1 U2694 ( .A(fifo_array[119]), .B(n4751), .Y(n281) );
  INVX1 U2695 ( .A(n281), .Y(n3131) );
  AND2X1 U2696 ( .A(fifo_array[107]), .B(n4751), .Y(n269) );
  INVX1 U2697 ( .A(n269), .Y(n3132) );
  AND2X1 U2698 ( .A(fifo_array[84]), .B(n4753), .Y(n244) );
  INVX1 U2699 ( .A(n244), .Y(n3133) );
  AND2X1 U2700 ( .A(fifo_array[72]), .B(n4753), .Y(n232) );
  INVX1 U2701 ( .A(n232), .Y(n3134) );
  AND2X1 U2702 ( .A(fifo_array[53]), .B(n4755), .Y(n211) );
  INVX1 U2703 ( .A(n211), .Y(n3135) );
  AND2X1 U2704 ( .A(fifo_array[41]), .B(n4755), .Y(n199) );
  INVX1 U2705 ( .A(n199), .Y(n3136) );
  AND2X1 U2706 ( .A(fifo_array[18]), .B(n4757), .Y(n173) );
  INVX1 U2707 ( .A(n173), .Y(n3137) );
  AND2X1 U2708 ( .A(fifo_array[6]), .B(n4756), .Y(n161) );
  INVX1 U2709 ( .A(n161), .Y(n3138) );
  AND2X1 U2710 ( .A(n3454), .B(n4758), .Y(n1355) );
  AND2X1 U2711 ( .A(n69), .B(n3457), .Y(n1290) );
  INVX1 U2712 ( .A(n1290), .Y(n3139) );
  AND2X1 U2713 ( .A(fifo_array[1063]), .B(n4695), .Y(n1261) );
  INVX1 U2714 ( .A(n1261), .Y(n3140) );
  AND2X1 U2715 ( .A(fifo_array[1054]), .B(n4694), .Y(n1252) );
  INVX1 U2716 ( .A(n1252), .Y(n3141) );
  AND2X1 U2717 ( .A(fifo_array[1033]), .B(n4697), .Y(n1230) );
  INVX1 U2718 ( .A(n1230), .Y(n3142) );
  AND2X1 U2719 ( .A(fifo_array[1021]), .B(n4696), .Y(n1218) );
  INVX1 U2720 ( .A(n1218), .Y(n3143) );
  AND2X1 U2721 ( .A(fifo_array[1004]), .B(n4699), .Y(n1200) );
  INVX1 U2722 ( .A(n1200), .Y(n3144) );
  AND2X1 U2723 ( .A(fifo_array[992]), .B(n4698), .Y(n1188) );
  INVX1 U2724 ( .A(n1188), .Y(n3145) );
  AND2X1 U2725 ( .A(fifo_array[971]), .B(n4701), .Y(n1166) );
  INVX1 U2726 ( .A(n1166), .Y(n3146) );
  AND2X1 U2727 ( .A(fifo_array[959]), .B(n4700), .Y(n1154) );
  INVX1 U2728 ( .A(n1154), .Y(n3147) );
  AND2X1 U2729 ( .A(fifo_array[934]), .B(n4703), .Y(n1128) );
  INVX1 U2730 ( .A(n1128), .Y(n3148) );
  AND2X1 U2731 ( .A(fifo_array[922]), .B(n4702), .Y(n1116) );
  INVX1 U2732 ( .A(n1116), .Y(n3149) );
  AND2X1 U2733 ( .A(fifo_array[901]), .B(n4705), .Y(n1094) );
  INVX1 U2734 ( .A(n1094), .Y(n3150) );
  AND2X1 U2735 ( .A(fifo_array[889]), .B(n4704), .Y(n1082) );
  INVX1 U2736 ( .A(n1082), .Y(n3151) );
  AND2X1 U2737 ( .A(fifo_array[871]), .B(n4706), .Y(n1063) );
  INVX1 U2738 ( .A(n1063), .Y(n3152) );
  AND2X1 U2739 ( .A(fifo_array[860]), .B(n4707), .Y(n1052) );
  INVX1 U2740 ( .A(n1052), .Y(n3153) );
  AND2X1 U2741 ( .A(fifo_array[841]), .B(n4709), .Y(n1031) );
  INVX1 U2742 ( .A(n1031), .Y(n3154) );
  AND2X1 U2743 ( .A(fifo_array[808]), .B(n4711), .Y(n997) );
  INVX1 U2744 ( .A(n997), .Y(n3155) );
  AND2X1 U2745 ( .A(fifo_array[771]), .B(n4713), .Y(n959) );
  INVX1 U2746 ( .A(n959), .Y(n3156) );
  AND2X1 U2747 ( .A(fifo_array[738]), .B(n4715), .Y(n925) );
  INVX1 U2748 ( .A(n925), .Y(n3157) );
  AND2X1 U2749 ( .A(fifo_array[694]), .B(n4717), .Y(n880) );
  INVX1 U2750 ( .A(n880), .Y(n3158) );
  AND2X1 U2751 ( .A(fifo_array[682]), .B(n4717), .Y(n868) );
  INVX1 U2752 ( .A(n868), .Y(n3159) );
  AND2X1 U2753 ( .A(fifo_array[661]), .B(n4719), .Y(n846) );
  INVX1 U2754 ( .A(n846), .Y(n3160) );
  AND2X1 U2755 ( .A(fifo_array[649]), .B(n4719), .Y(n834) );
  INVX1 U2756 ( .A(n834), .Y(n3161) );
  AND2X1 U2757 ( .A(fifo_array[621]), .B(n4721), .Y(n805) );
  INVX1 U2758 ( .A(n805), .Y(n3162) );
  AND2X1 U2759 ( .A(fifo_array[612]), .B(n4721), .Y(n796) );
  INVX1 U2760 ( .A(n796), .Y(n3163) );
  AND2X1 U2761 ( .A(fifo_array[591]), .B(n4723), .Y(n774) );
  INVX1 U2762 ( .A(n774), .Y(n3164) );
  AND2X1 U2763 ( .A(fifo_array[579]), .B(n4723), .Y(n762) );
  INVX1 U2764 ( .A(n762), .Y(n3165) );
  AND2X1 U2765 ( .A(fifo_array[562]), .B(n4725), .Y(n743) );
  INVX1 U2766 ( .A(n743), .Y(n3166) );
  AND2X1 U2767 ( .A(fifo_array[550]), .B(n4725), .Y(n731) );
  INVX1 U2768 ( .A(n731), .Y(n3167) );
  AND2X1 U2769 ( .A(fifo_array[529]), .B(n4727), .Y(n709) );
  INVX1 U2770 ( .A(n709), .Y(n3168) );
  AND2X1 U2771 ( .A(fifo_array[517]), .B(n4727), .Y(n697) );
  INVX1 U2772 ( .A(n697), .Y(n3169) );
  AND2X1 U2773 ( .A(fifo_array[492]), .B(n4729), .Y(n671) );
  INVX1 U2774 ( .A(n671), .Y(n3170) );
  AND2X1 U2775 ( .A(fifo_array[480]), .B(n4729), .Y(n659) );
  INVX1 U2776 ( .A(n659), .Y(n3171) );
  AND2X1 U2777 ( .A(fifo_array[459]), .B(n4731), .Y(n637) );
  INVX1 U2778 ( .A(n637), .Y(n3172) );
  AND2X1 U2779 ( .A(fifo_array[447]), .B(n4731), .Y(n625) );
  INVX1 U2780 ( .A(n625), .Y(n3173) );
  AND2X1 U2781 ( .A(fifo_array[429]), .B(n4732), .Y(n606) );
  INVX1 U2782 ( .A(n606), .Y(n3174) );
  AND2X1 U2783 ( .A(fifo_array[418]), .B(n4733), .Y(n595) );
  INVX1 U2784 ( .A(n595), .Y(n3175) );
  AND2X1 U2785 ( .A(fifo_array[399]), .B(n4735), .Y(n575) );
  INVX1 U2786 ( .A(n575), .Y(n3176) );
  AND2X1 U2787 ( .A(fifo_array[366]), .B(n4737), .Y(n541) );
  INVX1 U2788 ( .A(n541), .Y(n3177) );
  AND2X1 U2789 ( .A(fifo_array[329]), .B(n4739), .Y(n503) );
  INVX1 U2790 ( .A(n503), .Y(n3178) );
  AND2X1 U2791 ( .A(fifo_array[296]), .B(n4741), .Y(n468) );
  INVX1 U2792 ( .A(n468), .Y(n3179) );
  AND2X1 U2793 ( .A(fifo_array[252]), .B(n4743), .Y(n422) );
  INVX1 U2794 ( .A(n422), .Y(n3180) );
  AND2X1 U2795 ( .A(fifo_array[240]), .B(n4743), .Y(n410) );
  INVX1 U2796 ( .A(n410), .Y(n3181) );
  AND2X1 U2797 ( .A(fifo_array[219]), .B(n4745), .Y(n387) );
  INVX1 U2798 ( .A(n387), .Y(n3182) );
  AND2X1 U2799 ( .A(fifo_array[207]), .B(n4745), .Y(n375) );
  INVX1 U2800 ( .A(n375), .Y(n3183) );
  AND2X1 U2801 ( .A(fifo_array[179]), .B(n4747), .Y(n345) );
  INVX1 U2802 ( .A(n345), .Y(n3184) );
  AND2X1 U2803 ( .A(fifo_array[170]), .B(n4747), .Y(n336) );
  INVX1 U2804 ( .A(n336), .Y(n3185) );
  AND2X1 U2805 ( .A(fifo_array[149]), .B(n4749), .Y(n313) );
  INVX1 U2806 ( .A(n313), .Y(n3186) );
  AND2X1 U2807 ( .A(fifo_array[137]), .B(n4749), .Y(n301) );
  INVX1 U2808 ( .A(n301), .Y(n3187) );
  AND2X1 U2809 ( .A(fifo_array[120]), .B(n4751), .Y(n282) );
  INVX1 U2810 ( .A(n282), .Y(n3188) );
  AND2X1 U2811 ( .A(fifo_array[108]), .B(n4751), .Y(n270) );
  INVX1 U2812 ( .A(n270), .Y(n3189) );
  AND2X1 U2813 ( .A(fifo_array[87]), .B(n4753), .Y(n247) );
  INVX1 U2814 ( .A(n247), .Y(n3190) );
  AND2X1 U2815 ( .A(fifo_array[75]), .B(n4753), .Y(n235) );
  INVX1 U2816 ( .A(n235), .Y(n3191) );
  AND2X1 U2817 ( .A(fifo_array[50]), .B(n4755), .Y(n208) );
  INVX1 U2818 ( .A(n208), .Y(n3192) );
  AND2X1 U2819 ( .A(fifo_array[38]), .B(n4755), .Y(n196) );
  INVX1 U2820 ( .A(n196), .Y(n3193) );
  AND2X1 U2821 ( .A(fifo_array[17]), .B(n4757), .Y(n172) );
  INVX1 U2822 ( .A(n172), .Y(n3194) );
  AND2X1 U2823 ( .A(fifo_array[5]), .B(n4757), .Y(n160) );
  INVX1 U2824 ( .A(n160), .Y(n3195) );
  BUFX2 U2825 ( .A(n1300), .Y(n3196) );
  AND2X1 U2826 ( .A(n70), .B(n3457), .Y(n1289) );
  INVX1 U2827 ( .A(n1289), .Y(n3197) );
  AND2X1 U2828 ( .A(fifo_array[1067]), .B(n4695), .Y(n1265) );
  INVX1 U2829 ( .A(n1265), .Y(n3198) );
  AND2X1 U2830 ( .A(fifo_array[1055]), .B(n4694), .Y(n1253) );
  INVX1 U2831 ( .A(n1253), .Y(n3199) );
  AND2X1 U2832 ( .A(fifo_array[1029]), .B(n4697), .Y(n1226) );
  INVX1 U2833 ( .A(n1226), .Y(n3200) );
  AND2X1 U2834 ( .A(fifo_array[1020]), .B(n4696), .Y(n1217) );
  INVX1 U2835 ( .A(n1217), .Y(n3201) );
  AND2X1 U2836 ( .A(fifo_array[1005]), .B(n4699), .Y(n1201) );
  INVX1 U2837 ( .A(n1201), .Y(n3202) );
  AND2X1 U2838 ( .A(fifo_array[993]), .B(n4698), .Y(n1189) );
  INVX1 U2839 ( .A(n1189), .Y(n3203) );
  AND2X1 U2840 ( .A(fifo_array[970]), .B(n4701), .Y(n1165) );
  INVX1 U2841 ( .A(n1165), .Y(n3204) );
  AND2X1 U2842 ( .A(fifo_array[958]), .B(n4700), .Y(n1153) );
  INVX1 U2843 ( .A(n1153), .Y(n3205) );
  AND2X1 U2844 ( .A(fifo_array[935]), .B(n4703), .Y(n1129) );
  INVX1 U2845 ( .A(n1129), .Y(n3206) );
  AND2X1 U2846 ( .A(fifo_array[923]), .B(n4702), .Y(n1117) );
  INVX1 U2847 ( .A(n1117), .Y(n3207) );
  AND2X1 U2848 ( .A(fifo_array[900]), .B(n4705), .Y(n1093) );
  INVX1 U2849 ( .A(n1093), .Y(n3208) );
  AND2X1 U2850 ( .A(fifo_array[888]), .B(n4704), .Y(n1081) );
  INVX1 U2851 ( .A(n1081), .Y(n3209) );
  AND2X1 U2852 ( .A(fifo_array[870]), .B(n4706), .Y(n1062) );
  INVX1 U2853 ( .A(n1062), .Y(n3210) );
  AND2X1 U2854 ( .A(fifo_array[858]), .B(n4707), .Y(n1050) );
  INVX1 U2855 ( .A(n1050), .Y(n3211) );
  AND2X1 U2856 ( .A(fifo_array[842]), .B(n4709), .Y(n1032) );
  INVX1 U2857 ( .A(n1032), .Y(n3212) );
  AND2X1 U2858 ( .A(fifo_array[807]), .B(n4711), .Y(n996) );
  INVX1 U2859 ( .A(n996), .Y(n3213) );
  AND2X1 U2860 ( .A(fifo_array[772]), .B(n4713), .Y(n960) );
  INVX1 U2861 ( .A(n960), .Y(n3214) );
  AND2X1 U2862 ( .A(fifo_array[737]), .B(n4715), .Y(n924) );
  INVX1 U2863 ( .A(n924), .Y(n3215) );
  AND2X1 U2864 ( .A(fifo_array[695]), .B(n4717), .Y(n881) );
  INVX1 U2865 ( .A(n881), .Y(n3216) );
  AND2X1 U2866 ( .A(fifo_array[683]), .B(n4717), .Y(n869) );
  INVX1 U2867 ( .A(n869), .Y(n3217) );
  AND2X1 U2868 ( .A(fifo_array[660]), .B(n4719), .Y(n845) );
  INVX1 U2869 ( .A(n845), .Y(n3218) );
  AND2X1 U2870 ( .A(fifo_array[648]), .B(n4719), .Y(n833) );
  INVX1 U2871 ( .A(n833), .Y(n3219) );
  AND2X1 U2872 ( .A(fifo_array[625]), .B(n4721), .Y(n809) );
  INVX1 U2873 ( .A(n809), .Y(n3220) );
  AND2X1 U2874 ( .A(fifo_array[613]), .B(n4721), .Y(n797) );
  INVX1 U2875 ( .A(n797), .Y(n3221) );
  AND2X1 U2876 ( .A(fifo_array[587]), .B(n4723), .Y(n770) );
  INVX1 U2877 ( .A(n770), .Y(n3222) );
  AND2X1 U2878 ( .A(fifo_array[578]), .B(n4723), .Y(n761) );
  INVX1 U2879 ( .A(n761), .Y(n3223) );
  AND2X1 U2880 ( .A(fifo_array[563]), .B(n4725), .Y(n744) );
  INVX1 U2881 ( .A(n744), .Y(n3224) );
  AND2X1 U2882 ( .A(fifo_array[551]), .B(n4725), .Y(n732) );
  INVX1 U2883 ( .A(n732), .Y(n3225) );
  AND2X1 U2884 ( .A(fifo_array[528]), .B(n4727), .Y(n708) );
  INVX1 U2885 ( .A(n708), .Y(n3226) );
  AND2X1 U2886 ( .A(fifo_array[516]), .B(n4727), .Y(n696) );
  INVX1 U2887 ( .A(n696), .Y(n3227) );
  AND2X1 U2888 ( .A(fifo_array[493]), .B(n4729), .Y(n672) );
  INVX1 U2889 ( .A(n672), .Y(n3228) );
  AND2X1 U2890 ( .A(fifo_array[481]), .B(n4729), .Y(n660) );
  INVX1 U2891 ( .A(n660), .Y(n3229) );
  AND2X1 U2892 ( .A(fifo_array[458]), .B(n4731), .Y(n636) );
  INVX1 U2893 ( .A(n636), .Y(n3230) );
  AND2X1 U2894 ( .A(fifo_array[446]), .B(n4731), .Y(n624) );
  INVX1 U2895 ( .A(n624), .Y(n3231) );
  AND2X1 U2896 ( .A(fifo_array[428]), .B(n4732), .Y(n605) );
  INVX1 U2897 ( .A(n605), .Y(n3232) );
  AND2X1 U2898 ( .A(fifo_array[416]), .B(n4732), .Y(n593) );
  INVX1 U2899 ( .A(n593), .Y(n3233) );
  AND2X1 U2900 ( .A(fifo_array[400]), .B(n4735), .Y(n576) );
  INVX1 U2901 ( .A(n576), .Y(n3234) );
  AND2X1 U2902 ( .A(fifo_array[365]), .B(n4737), .Y(n540) );
  INVX1 U2903 ( .A(n540), .Y(n3235) );
  AND2X1 U2904 ( .A(fifo_array[330]), .B(n4739), .Y(n504) );
  INVX1 U2905 ( .A(n504), .Y(n3236) );
  AND2X1 U2906 ( .A(fifo_array[295]), .B(n4741), .Y(n467) );
  INVX1 U2907 ( .A(n467), .Y(n3237) );
  AND2X1 U2908 ( .A(fifo_array[253]), .B(n4743), .Y(n423) );
  INVX1 U2909 ( .A(n423), .Y(n3238) );
  AND2X1 U2910 ( .A(fifo_array[241]), .B(n4743), .Y(n411) );
  INVX1 U2911 ( .A(n411), .Y(n3239) );
  AND2X1 U2912 ( .A(fifo_array[218]), .B(n4745), .Y(n386) );
  INVX1 U2913 ( .A(n386), .Y(n3240) );
  AND2X1 U2914 ( .A(fifo_array[206]), .B(n4745), .Y(n374) );
  INVX1 U2915 ( .A(n374), .Y(n3241) );
  AND2X1 U2916 ( .A(fifo_array[183]), .B(n4747), .Y(n349) );
  INVX1 U2917 ( .A(n349), .Y(n3242) );
  AND2X1 U2918 ( .A(fifo_array[171]), .B(n4747), .Y(n337) );
  INVX1 U2919 ( .A(n337), .Y(n3243) );
  AND2X1 U2920 ( .A(fifo_array[145]), .B(n4749), .Y(n309) );
  INVX1 U2921 ( .A(n309), .Y(n3244) );
  AND2X1 U2922 ( .A(fifo_array[136]), .B(n4749), .Y(n300) );
  INVX1 U2923 ( .A(n300), .Y(n3245) );
  AND2X1 U2924 ( .A(fifo_array[121]), .B(n4751), .Y(n283) );
  INVX1 U2925 ( .A(n283), .Y(n3246) );
  AND2X1 U2926 ( .A(fifo_array[109]), .B(n4751), .Y(n271) );
  INVX1 U2927 ( .A(n271), .Y(n3247) );
  AND2X1 U2928 ( .A(fifo_array[86]), .B(n4753), .Y(n246) );
  INVX1 U2929 ( .A(n246), .Y(n3248) );
  AND2X1 U2930 ( .A(fifo_array[74]), .B(n4753), .Y(n234) );
  INVX1 U2931 ( .A(n234), .Y(n3249) );
  AND2X1 U2932 ( .A(fifo_array[51]), .B(n4755), .Y(n209) );
  INVX1 U2933 ( .A(n209), .Y(n3250) );
  AND2X1 U2934 ( .A(fifo_array[39]), .B(n4755), .Y(n197) );
  INVX1 U2935 ( .A(n197), .Y(n3251) );
  AND2X1 U2936 ( .A(fifo_array[16]), .B(n4757), .Y(n171) );
  INVX1 U2937 ( .A(n171), .Y(n3252) );
  AND2X1 U2938 ( .A(fifo_array[4]), .B(n4757), .Y(n159) );
  INVX1 U2939 ( .A(n159), .Y(n3253) );
  BUFX2 U2940 ( .A(n1299), .Y(n3254) );
  BUFX2 U2941 ( .A(n1345), .Y(n3255) );
  INVX1 U2942 ( .A(n1357), .Y(n3256) );
  BUFX2 U2943 ( .A(n1356), .Y(n3257) );
  BUFX2 U2944 ( .A(n1358), .Y(n3258) );
  AND2X1 U2945 ( .A(n71), .B(n3457), .Y(n1287) );
  INVX1 U2946 ( .A(n1287), .Y(n3259) );
  AND2X1 U2947 ( .A(fifo_array[1072]), .B(n4695), .Y(n1270) );
  INVX1 U2948 ( .A(n1270), .Y(n3260) );
  AND2X1 U2949 ( .A(fifo_array[1060]), .B(n4695), .Y(n1258) );
  INVX1 U2950 ( .A(n1258), .Y(n3261) );
  AND2X1 U2951 ( .A(fifo_array[1039]), .B(n4697), .Y(n1236) );
  INVX1 U2952 ( .A(n1236), .Y(n3262) );
  AND2X1 U2953 ( .A(fifo_array[1027]), .B(n4697), .Y(n1224) );
  INVX1 U2954 ( .A(n1224), .Y(n3263) );
  AND2X1 U2955 ( .A(fifo_array[995]), .B(n4699), .Y(n1191) );
  INVX1 U2956 ( .A(n1191), .Y(n3264) );
  AND2X1 U2957 ( .A(fifo_array[986]), .B(n4699), .Y(n1182) );
  INVX1 U2958 ( .A(n1182), .Y(n3265) );
  AND2X1 U2959 ( .A(fifo_array[965]), .B(n4701), .Y(n1160) );
  INVX1 U2960 ( .A(n1160), .Y(n3266) );
  AND2X1 U2961 ( .A(fifo_array[953]), .B(n4701), .Y(n1148) );
  INVX1 U2962 ( .A(n1148), .Y(n3267) );
  AND2X1 U2963 ( .A(fifo_array[932]), .B(n4703), .Y(n1126) );
  INVX1 U2964 ( .A(n1126), .Y(n3268) );
  AND2X1 U2965 ( .A(fifo_array[920]), .B(n4703), .Y(n1114) );
  INVX1 U2966 ( .A(n1114), .Y(n3269) );
  AND2X1 U2967 ( .A(fifo_array[899]), .B(n4705), .Y(n1092) );
  INVX1 U2968 ( .A(n1092), .Y(n3270) );
  AND2X1 U2969 ( .A(fifo_array[887]), .B(n4705), .Y(n1080) );
  INVX1 U2970 ( .A(n1080), .Y(n3271) );
  AND2X1 U2971 ( .A(fifo_array[876]), .B(n4707), .Y(n1068) );
  INVX1 U2972 ( .A(n1068), .Y(n3272) );
  AND2X1 U2973 ( .A(fifo_array[836]), .B(n4708), .Y(n1026) );
  INVX1 U2974 ( .A(n1026), .Y(n3273) );
  AND2X1 U2975 ( .A(fifo_array[824]), .B(n4709), .Y(n1014) );
  INVX1 U2976 ( .A(n1014), .Y(n3274) );
  AND2X1 U2977 ( .A(fifo_array[803]), .B(n4710), .Y(n992) );
  INVX1 U2978 ( .A(n992), .Y(n3275) );
  AND2X1 U2979 ( .A(fifo_array[792]), .B(n4711), .Y(n981) );
  INVX1 U2980 ( .A(n981), .Y(n3276) );
  AND2X1 U2981 ( .A(fifo_array[770]), .B(n4712), .Y(n958) );
  INVX1 U2982 ( .A(n958), .Y(n3277) );
  AND2X1 U2983 ( .A(fifo_array[759]), .B(n4713), .Y(n947) );
  INVX1 U2984 ( .A(n947), .Y(n3278) );
  AND2X1 U2985 ( .A(fifo_array[743]), .B(n4714), .Y(n930) );
  INVX1 U2986 ( .A(n930), .Y(n3279) );
  AND2X1 U2987 ( .A(fifo_array[726]), .B(n4715), .Y(n913) );
  INVX1 U2988 ( .A(n913), .Y(n3280) );
  AND2X1 U2989 ( .A(fifo_array[696]), .B(n4717), .Y(n882) );
  INVX1 U2990 ( .A(n882), .Y(n3281) );
  AND2X1 U2991 ( .A(fifo_array[684]), .B(n4717), .Y(n870) );
  INVX1 U2992 ( .A(n870), .Y(n3282) );
  AND2X1 U2993 ( .A(fifo_array[663]), .B(n4719), .Y(n848) );
  INVX1 U2994 ( .A(n848), .Y(n3283) );
  AND2X1 U2995 ( .A(fifo_array[651]), .B(n4719), .Y(n836) );
  INVX1 U2996 ( .A(n836), .Y(n3284) );
  AND2X1 U2997 ( .A(fifo_array[630]), .B(n4721), .Y(n814) );
  INVX1 U2998 ( .A(n814), .Y(n3285) );
  AND2X1 U2999 ( .A(fifo_array[618]), .B(n4721), .Y(n802) );
  INVX1 U3000 ( .A(n802), .Y(n3286) );
  AND2X1 U3001 ( .A(fifo_array[597]), .B(n4723), .Y(n780) );
  INVX1 U3002 ( .A(n780), .Y(n3287) );
  AND2X1 U3003 ( .A(fifo_array[585]), .B(n4723), .Y(n768) );
  INVX1 U3004 ( .A(n768), .Y(n3288) );
  AND2X1 U3005 ( .A(fifo_array[553]), .B(n4725), .Y(n734) );
  INVX1 U3006 ( .A(n734), .Y(n3289) );
  AND2X1 U3007 ( .A(fifo_array[544]), .B(n4725), .Y(n725) );
  INVX1 U3008 ( .A(n725), .Y(n3290) );
  AND2X1 U3009 ( .A(fifo_array[523]), .B(n4727), .Y(n703) );
  INVX1 U3010 ( .A(n703), .Y(n3291) );
  AND2X1 U3011 ( .A(fifo_array[511]), .B(n4727), .Y(n691) );
  INVX1 U3012 ( .A(n691), .Y(n3292) );
  AND2X1 U3013 ( .A(fifo_array[490]), .B(n4729), .Y(n669) );
  INVX1 U3014 ( .A(n669), .Y(n3293) );
  AND2X1 U3015 ( .A(fifo_array[478]), .B(n4729), .Y(n657) );
  INVX1 U3016 ( .A(n657), .Y(n3294) );
  AND2X1 U3017 ( .A(fifo_array[457]), .B(n4731), .Y(n635) );
  INVX1 U3018 ( .A(n635), .Y(n3295) );
  AND2X1 U3019 ( .A(fifo_array[445]), .B(n4731), .Y(n623) );
  INVX1 U3020 ( .A(n623), .Y(n3296) );
  AND2X1 U3021 ( .A(fifo_array[434]), .B(n4733), .Y(n611) );
  INVX1 U3022 ( .A(n611), .Y(n3297) );
  AND2X1 U3023 ( .A(fifo_array[394]), .B(n4734), .Y(n570) );
  INVX1 U3024 ( .A(n570), .Y(n3298) );
  AND2X1 U3025 ( .A(fifo_array[382]), .B(n4734), .Y(n558) );
  INVX1 U3026 ( .A(n558), .Y(n3299) );
  AND2X1 U3027 ( .A(fifo_array[361]), .B(n4736), .Y(n536) );
  INVX1 U3028 ( .A(n536), .Y(n3300) );
  AND2X1 U3029 ( .A(fifo_array[350]), .B(n4737), .Y(n525) );
  INVX1 U3030 ( .A(n525), .Y(n3301) );
  AND2X1 U3031 ( .A(fifo_array[328]), .B(n4738), .Y(n502) );
  INVX1 U3032 ( .A(n502), .Y(n3302) );
  AND2X1 U3033 ( .A(fifo_array[317]), .B(n4739), .Y(n491) );
  INVX1 U3034 ( .A(n491), .Y(n3303) );
  AND2X1 U3035 ( .A(fifo_array[301]), .B(n4740), .Y(n473) );
  INVX1 U3036 ( .A(n473), .Y(n3304) );
  AND2X1 U3037 ( .A(fifo_array[284]), .B(n4741), .Y(n456) );
  INVX1 U3038 ( .A(n456), .Y(n3305) );
  AND2X1 U3039 ( .A(fifo_array[254]), .B(n4743), .Y(n424) );
  INVX1 U3040 ( .A(n424), .Y(n3306) );
  AND2X1 U3041 ( .A(fifo_array[242]), .B(n4743), .Y(n412) );
  INVX1 U3042 ( .A(n412), .Y(n3307) );
  AND2X1 U3043 ( .A(fifo_array[221]), .B(n4745), .Y(n389) );
  INVX1 U3044 ( .A(n389), .Y(n3308) );
  AND2X1 U3045 ( .A(fifo_array[209]), .B(n4745), .Y(n377) );
  INVX1 U3046 ( .A(n377), .Y(n3309) );
  AND2X1 U3047 ( .A(fifo_array[188]), .B(n4747), .Y(n354) );
  INVX1 U3048 ( .A(n354), .Y(n3310) );
  AND2X1 U3049 ( .A(fifo_array[176]), .B(n4747), .Y(n342) );
  INVX1 U3050 ( .A(n342), .Y(n3311) );
  AND2X1 U3051 ( .A(fifo_array[155]), .B(n4749), .Y(n319) );
  INVX1 U3052 ( .A(n319), .Y(n3312) );
  AND2X1 U3053 ( .A(fifo_array[143]), .B(n4749), .Y(n307) );
  INVX1 U3054 ( .A(n307), .Y(n3313) );
  AND2X1 U3055 ( .A(fifo_array[111]), .B(n4751), .Y(n273) );
  INVX1 U3056 ( .A(n273), .Y(n3314) );
  AND2X1 U3057 ( .A(fifo_array[102]), .B(n4751), .Y(n264) );
  INVX1 U3058 ( .A(n264), .Y(n3315) );
  AND2X1 U3059 ( .A(fifo_array[81]), .B(n4753), .Y(n241) );
  INVX1 U3060 ( .A(n241), .Y(n3316) );
  AND2X1 U3061 ( .A(fifo_array[69]), .B(n4753), .Y(n229) );
  INVX1 U3062 ( .A(n229), .Y(n3317) );
  AND2X1 U3063 ( .A(fifo_array[48]), .B(n4755), .Y(n206) );
  INVX1 U3064 ( .A(n206), .Y(n3318) );
  AND2X1 U3065 ( .A(fifo_array[36]), .B(n4755), .Y(n194) );
  INVX1 U3066 ( .A(n194), .Y(n3319) );
  AND2X1 U3067 ( .A(fifo_array[15]), .B(n4757), .Y(n170) );
  INVX1 U3068 ( .A(n170), .Y(n3320) );
  AND2X1 U3069 ( .A(fifo_array[3]), .B(n4757), .Y(n158) );
  INVX1 U3070 ( .A(n158), .Y(n3321) );
  BUFX2 U3071 ( .A(n1301), .Y(n3322) );
  INVX1 U3072 ( .A(n1347), .Y(n3323) );
  BUFX2 U3073 ( .A(n1346), .Y(n3324) );
  BUFX2 U3074 ( .A(n1349), .Y(n3325) );
  AND2X1 U3075 ( .A(fifo_array[1073]), .B(n4695), .Y(n1271) );
  INVX1 U3076 ( .A(n1271), .Y(n3326) );
  AND2X1 U3077 ( .A(fifo_array[1061]), .B(n4694), .Y(n1259) );
  INVX1 U3078 ( .A(n1259), .Y(n3327) );
  AND2X1 U3079 ( .A(fifo_array[1038]), .B(n4697), .Y(n1235) );
  INVX1 U3080 ( .A(n1235), .Y(n3328) );
  AND2X1 U3081 ( .A(fifo_array[1026]), .B(n4696), .Y(n1223) );
  INVX1 U3082 ( .A(n1223), .Y(n3329) );
  AND2X1 U3083 ( .A(fifo_array[999]), .B(n4699), .Y(n1195) );
  INVX1 U3084 ( .A(n1195), .Y(n3330) );
  AND2X1 U3085 ( .A(fifo_array[987]), .B(n4698), .Y(n1183) );
  INVX1 U3086 ( .A(n1183), .Y(n3331) );
  AND2X1 U3087 ( .A(fifo_array[961]), .B(n4701), .Y(n1156) );
  INVX1 U3088 ( .A(n1156), .Y(n3332) );
  AND2X1 U3089 ( .A(fifo_array[952]), .B(n4700), .Y(n1147) );
  INVX1 U3090 ( .A(n1147), .Y(n3333) );
  AND2X1 U3091 ( .A(fifo_array[933]), .B(n4703), .Y(n1127) );
  INVX1 U3092 ( .A(n1127), .Y(n3334) );
  AND2X1 U3093 ( .A(fifo_array[921]), .B(n4702), .Y(n1115) );
  INVX1 U3094 ( .A(n1115), .Y(n3335) );
  AND2X1 U3095 ( .A(fifo_array[898]), .B(n4705), .Y(n1091) );
  INVX1 U3096 ( .A(n1091), .Y(n3336) );
  AND2X1 U3097 ( .A(fifo_array[886]), .B(n4704), .Y(n1079) );
  INVX1 U3098 ( .A(n1079), .Y(n3337) );
  AND2X1 U3099 ( .A(fifo_array[875]), .B(n4707), .Y(n1067) );
  INVX1 U3100 ( .A(n1067), .Y(n3338) );
  AND2X1 U3101 ( .A(fifo_array[837]), .B(n4708), .Y(n1027) );
  INVX1 U3102 ( .A(n1027), .Y(n3339) );
  AND2X1 U3103 ( .A(fifo_array[826]), .B(n4709), .Y(n1016) );
  INVX1 U3104 ( .A(n1016), .Y(n3340) );
  AND2X1 U3105 ( .A(fifo_array[802]), .B(n4710), .Y(n991) );
  INVX1 U3106 ( .A(n991), .Y(n3341) );
  AND2X1 U3107 ( .A(fifo_array[790]), .B(n4710), .Y(n979) );
  INVX1 U3108 ( .A(n979), .Y(n3342) );
  AND2X1 U3109 ( .A(fifo_array[777]), .B(n4712), .Y(n965) );
  INVX1 U3110 ( .A(n965), .Y(n3343) );
  AND2X1 U3111 ( .A(fifo_array[760]), .B(n4713), .Y(n948) );
  INVX1 U3112 ( .A(n948), .Y(n3344) );
  AND2X1 U3113 ( .A(fifo_array[736]), .B(n4714), .Y(n923) );
  INVX1 U3114 ( .A(n923), .Y(n3345) );
  AND2X1 U3115 ( .A(fifo_array[725]), .B(n4715), .Y(n912) );
  INVX1 U3116 ( .A(n912), .Y(n3346) );
  AND2X1 U3117 ( .A(fifo_array[697]), .B(n4717), .Y(n883) );
  INVX1 U3118 ( .A(n883), .Y(n3347) );
  AND2X1 U3119 ( .A(fifo_array[685]), .B(n4717), .Y(n871) );
  INVX1 U3120 ( .A(n871), .Y(n3348) );
  AND2X1 U3121 ( .A(fifo_array[662]), .B(n4719), .Y(n847) );
  INVX1 U3122 ( .A(n847), .Y(n3349) );
  AND2X1 U3123 ( .A(fifo_array[650]), .B(n4719), .Y(n835) );
  INVX1 U3124 ( .A(n835), .Y(n3350) );
  AND2X1 U3125 ( .A(fifo_array[631]), .B(n4721), .Y(n815) );
  INVX1 U3126 ( .A(n815), .Y(n3351) );
  AND2X1 U3127 ( .A(fifo_array[619]), .B(n4721), .Y(n803) );
  INVX1 U3128 ( .A(n803), .Y(n3352) );
  AND2X1 U3129 ( .A(fifo_array[596]), .B(n4723), .Y(n779) );
  INVX1 U3130 ( .A(n779), .Y(n3353) );
  AND2X1 U3131 ( .A(fifo_array[584]), .B(n4723), .Y(n767) );
  INVX1 U3132 ( .A(n767), .Y(n3354) );
  AND2X1 U3133 ( .A(fifo_array[557]), .B(n4725), .Y(n738) );
  INVX1 U3134 ( .A(n738), .Y(n3355) );
  AND2X1 U3135 ( .A(fifo_array[545]), .B(n4725), .Y(n726) );
  INVX1 U3136 ( .A(n726), .Y(n3356) );
  AND2X1 U3137 ( .A(fifo_array[519]), .B(n4727), .Y(n699) );
  INVX1 U3138 ( .A(n699), .Y(n3357) );
  AND2X1 U3139 ( .A(fifo_array[510]), .B(n4727), .Y(n690) );
  INVX1 U3140 ( .A(n690), .Y(n3358) );
  AND2X1 U3141 ( .A(fifo_array[491]), .B(n4729), .Y(n670) );
  INVX1 U3142 ( .A(n670), .Y(n3359) );
  AND2X1 U3143 ( .A(fifo_array[479]), .B(n4729), .Y(n658) );
  INVX1 U3144 ( .A(n658), .Y(n3360) );
  AND2X1 U3145 ( .A(fifo_array[456]), .B(n4731), .Y(n634) );
  INVX1 U3146 ( .A(n634), .Y(n3361) );
  AND2X1 U3147 ( .A(fifo_array[444]), .B(n4731), .Y(n622) );
  INVX1 U3148 ( .A(n622), .Y(n3362) );
  AND2X1 U3149 ( .A(fifo_array[433]), .B(n4733), .Y(n610) );
  INVX1 U3150 ( .A(n610), .Y(n3363) );
  AND2X1 U3151 ( .A(fifo_array[395]), .B(n4734), .Y(n571) );
  INVX1 U3152 ( .A(n571), .Y(n3364) );
  AND2X1 U3153 ( .A(fifo_array[384]), .B(n4735), .Y(n560) );
  INVX1 U3154 ( .A(n560), .Y(n3365) );
  AND2X1 U3155 ( .A(fifo_array[360]), .B(n4736), .Y(n535) );
  INVX1 U3156 ( .A(n535), .Y(n3366) );
  AND2X1 U3157 ( .A(fifo_array[348]), .B(n4736), .Y(n523) );
  INVX1 U3158 ( .A(n523), .Y(n3367) );
  AND2X1 U3159 ( .A(fifo_array[335]), .B(n4738), .Y(n509) );
  INVX1 U3160 ( .A(n509), .Y(n3368) );
  AND2X1 U3161 ( .A(fifo_array[318]), .B(n4739), .Y(n492) );
  INVX1 U3162 ( .A(n492), .Y(n3369) );
  AND2X1 U3163 ( .A(fifo_array[294]), .B(n4740), .Y(n466) );
  INVX1 U3164 ( .A(n466), .Y(n3370) );
  AND2X1 U3165 ( .A(fifo_array[283]), .B(n4741), .Y(n455) );
  INVX1 U3166 ( .A(n455), .Y(n3371) );
  AND2X1 U3167 ( .A(fifo_array[255]), .B(n4743), .Y(n425) );
  INVX1 U3168 ( .A(n425), .Y(n3372) );
  AND2X1 U3169 ( .A(fifo_array[243]), .B(n4742), .Y(n413) );
  INVX1 U3170 ( .A(n413), .Y(n3373) );
  AND2X1 U3171 ( .A(fifo_array[220]), .B(n4745), .Y(n388) );
  INVX1 U3172 ( .A(n388), .Y(n3374) );
  AND2X1 U3173 ( .A(fifo_array[208]), .B(n4744), .Y(n376) );
  INVX1 U3174 ( .A(n376), .Y(n3375) );
  AND2X1 U3175 ( .A(fifo_array[189]), .B(n4747), .Y(n355) );
  INVX1 U3176 ( .A(n355), .Y(n3376) );
  AND2X1 U3177 ( .A(fifo_array[177]), .B(n4746), .Y(n343) );
  INVX1 U3178 ( .A(n343), .Y(n3377) );
  AND2X1 U3179 ( .A(fifo_array[154]), .B(n4749), .Y(n318) );
  INVX1 U3180 ( .A(n318), .Y(n3378) );
  AND2X1 U3181 ( .A(fifo_array[142]), .B(n4748), .Y(n306) );
  INVX1 U3182 ( .A(n306), .Y(n3379) );
  AND2X1 U3183 ( .A(fifo_array[115]), .B(n4751), .Y(n277) );
  INVX1 U3184 ( .A(n277), .Y(n3380) );
  AND2X1 U3185 ( .A(fifo_array[103]), .B(n4750), .Y(n265) );
  INVX1 U3186 ( .A(n265), .Y(n3381) );
  AND2X1 U3187 ( .A(fifo_array[77]), .B(n4753), .Y(n237) );
  INVX1 U3188 ( .A(n237), .Y(n3382) );
  AND2X1 U3189 ( .A(fifo_array[68]), .B(n4752), .Y(n228) );
  INVX1 U3190 ( .A(n228), .Y(n3383) );
  AND2X1 U3191 ( .A(fifo_array[49]), .B(n4755), .Y(n207) );
  INVX1 U3192 ( .A(n207), .Y(n3384) );
  AND2X1 U3193 ( .A(fifo_array[37]), .B(n4754), .Y(n195) );
  INVX1 U3194 ( .A(n195), .Y(n3385) );
  AND2X1 U3195 ( .A(fifo_array[14]), .B(n4757), .Y(n169) );
  INVX1 U3196 ( .A(n169), .Y(n3386) );
  AND2X1 U3197 ( .A(fifo_array[2]), .B(n4756), .Y(n157) );
  INVX1 U3198 ( .A(n157), .Y(n3387) );
  BUFX2 U3199 ( .A(n1353), .Y(n3388) );
  OR2X1 U3200 ( .A(n95), .B(n4814), .Y(n1360) );
  INVX1 U3201 ( .A(n1360), .Y(n3389) );
  INVX1 U3202 ( .A(n1293), .Y(n3390) );
  AND2X1 U3203 ( .A(fifo_array[1070]), .B(n4695), .Y(n1268) );
  INVX1 U3204 ( .A(n1268), .Y(n3391) );
  AND2X1 U3205 ( .A(fifo_array[1058]), .B(n4695), .Y(n1256) );
  INVX1 U3206 ( .A(n1256), .Y(n3392) );
  AND2X1 U3207 ( .A(fifo_array[1037]), .B(n4697), .Y(n1234) );
  INVX1 U3208 ( .A(n1234), .Y(n3393) );
  AND2X1 U3209 ( .A(fifo_array[1025]), .B(n4697), .Y(n1222) );
  INVX1 U3210 ( .A(n1222), .Y(n3394) );
  AND2X1 U3211 ( .A(fifo_array[1000]), .B(n4699), .Y(n1196) );
  INVX1 U3212 ( .A(n1196), .Y(n3395) );
  AND2X1 U3213 ( .A(fifo_array[988]), .B(n4699), .Y(n1184) );
  INVX1 U3214 ( .A(n1184), .Y(n3396) );
  AND2X1 U3215 ( .A(fifo_array[967]), .B(n4701), .Y(n1162) );
  INVX1 U3216 ( .A(n1162), .Y(n3397) );
  AND2X1 U3217 ( .A(fifo_array[955]), .B(n4701), .Y(n1150) );
  INVX1 U3218 ( .A(n1150), .Y(n3398) );
  AND2X1 U3219 ( .A(fifo_array[927]), .B(n4703), .Y(n1121) );
  INVX1 U3220 ( .A(n1121), .Y(n3399) );
  AND2X1 U3221 ( .A(fifo_array[918]), .B(n4703), .Y(n1112) );
  INVX1 U3222 ( .A(n1112), .Y(n3400) );
  AND2X1 U3223 ( .A(fifo_array[897]), .B(n4705), .Y(n1090) );
  INVX1 U3224 ( .A(n1090), .Y(n3401) );
  AND2X1 U3225 ( .A(fifo_array[885]), .B(n4705), .Y(n1078) );
  INVX1 U3226 ( .A(n1078), .Y(n3402) );
  AND2X1 U3227 ( .A(fifo_array[874]), .B(n4707), .Y(n1066) );
  INVX1 U3228 ( .A(n1066), .Y(n3403) );
  AND2X1 U3229 ( .A(fifo_array[838]), .B(n4708), .Y(n1028) );
  INVX1 U3230 ( .A(n1028), .Y(n3404) );
  AND2X1 U3231 ( .A(fifo_array[827]), .B(n4709), .Y(n1017) );
  INVX1 U3232 ( .A(n1017), .Y(n3405) );
  AND2X1 U3233 ( .A(fifo_array[811]), .B(n4710), .Y(n1000) );
  INVX1 U3234 ( .A(n1000), .Y(n3406) );
  AND2X1 U3235 ( .A(fifo_array[794]), .B(n4711), .Y(n983) );
  INVX1 U3236 ( .A(n983), .Y(n3407) );
  AND2X1 U3237 ( .A(fifo_array[768]), .B(n4712), .Y(n956) );
  INVX1 U3238 ( .A(n956), .Y(n3408) );
  AND2X1 U3239 ( .A(fifo_array[756]), .B(n4712), .Y(n944) );
  INVX1 U3240 ( .A(n944), .Y(n3409) );
  AND2X1 U3241 ( .A(fifo_array[735]), .B(n4714), .Y(n922) );
  INVX1 U3242 ( .A(n922), .Y(n3410) );
  AND2X1 U3243 ( .A(fifo_array[724]), .B(n4715), .Y(n911) );
  INVX1 U3244 ( .A(n911), .Y(n3411) );
  AND2X1 U3245 ( .A(fifo_array[698]), .B(n4717), .Y(n884) );
  INVX1 U3246 ( .A(n884), .Y(n3412) );
  AND2X1 U3247 ( .A(fifo_array[686]), .B(n4716), .Y(n872) );
  INVX1 U3248 ( .A(n872), .Y(n3413) );
  AND2X1 U3249 ( .A(fifo_array[665]), .B(n4719), .Y(n850) );
  INVX1 U3250 ( .A(n850), .Y(n3414) );
  AND2X1 U3251 ( .A(fifo_array[653]), .B(n4718), .Y(n838) );
  INVX1 U3252 ( .A(n838), .Y(n3415) );
  AND2X1 U3253 ( .A(fifo_array[628]), .B(n4721), .Y(n812) );
  INVX1 U3254 ( .A(n812), .Y(n3416) );
  AND2X1 U3255 ( .A(fifo_array[616]), .B(n4720), .Y(n800) );
  INVX1 U3256 ( .A(n800), .Y(n3417) );
  AND2X1 U3257 ( .A(fifo_array[595]), .B(n4723), .Y(n778) );
  INVX1 U3258 ( .A(n778), .Y(n3418) );
  AND2X1 U3259 ( .A(fifo_array[583]), .B(n4722), .Y(n766) );
  INVX1 U3260 ( .A(n766), .Y(n3419) );
  AND2X1 U3261 ( .A(fifo_array[558]), .B(n4725), .Y(n739) );
  INVX1 U3262 ( .A(n739), .Y(n3420) );
  AND2X1 U3263 ( .A(fifo_array[546]), .B(n4724), .Y(n727) );
  INVX1 U3264 ( .A(n727), .Y(n3421) );
  AND2X1 U3265 ( .A(fifo_array[525]), .B(n4727), .Y(n705) );
  INVX1 U3266 ( .A(n705), .Y(n3422) );
  AND2X1 U3267 ( .A(fifo_array[513]), .B(n4726), .Y(n693) );
  INVX1 U3268 ( .A(n693), .Y(n3423) );
  AND2X1 U3269 ( .A(fifo_array[485]), .B(n4729), .Y(n664) );
  INVX1 U3270 ( .A(n664), .Y(n3424) );
  AND2X1 U3271 ( .A(fifo_array[476]), .B(n4728), .Y(n655) );
  INVX1 U3272 ( .A(n655), .Y(n3425) );
  AND2X1 U3273 ( .A(fifo_array[455]), .B(n4731), .Y(n633) );
  INVX1 U3274 ( .A(n633), .Y(n3426) );
  AND2X1 U3275 ( .A(fifo_array[443]), .B(n4730), .Y(n621) );
  INVX1 U3276 ( .A(n621), .Y(n3427) );
  AND2X1 U3277 ( .A(fifo_array[432]), .B(n4733), .Y(n609) );
  INVX1 U3278 ( .A(n609), .Y(n3428) );
  AND2X1 U3279 ( .A(fifo_array[396]), .B(n4734), .Y(n572) );
  INVX1 U3280 ( .A(n572), .Y(n3429) );
  AND2X1 U3281 ( .A(fifo_array[385]), .B(n4735), .Y(n561) );
  INVX1 U3282 ( .A(n561), .Y(n3430) );
  AND2X1 U3283 ( .A(fifo_array[369]), .B(n4736), .Y(n544) );
  INVX1 U3284 ( .A(n544), .Y(n3431) );
  AND2X1 U3285 ( .A(fifo_array[352]), .B(n4737), .Y(n527) );
  INVX1 U3286 ( .A(n527), .Y(n3432) );
  AND2X1 U3287 ( .A(fifo_array[326]), .B(n4738), .Y(n500) );
  INVX1 U3288 ( .A(n500), .Y(n3433) );
  AND2X1 U3289 ( .A(fifo_array[314]), .B(n4738), .Y(n488) );
  INVX1 U3290 ( .A(n488), .Y(n3434) );
  AND2X1 U3291 ( .A(fifo_array[293]), .B(n4740), .Y(n465) );
  INVX1 U3292 ( .A(n465), .Y(n3435) );
  AND2X1 U3293 ( .A(fifo_array[282]), .B(n4741), .Y(n454) );
  INVX1 U3294 ( .A(n454), .Y(n3436) );
  AND2X1 U3295 ( .A(fifo_array[256]), .B(n4743), .Y(n426) );
  INVX1 U3296 ( .A(n426), .Y(n3437) );
  AND2X1 U3297 ( .A(fifo_array[244]), .B(n4743), .Y(n414) );
  INVX1 U3298 ( .A(n414), .Y(n3438) );
  AND2X1 U3299 ( .A(fifo_array[223]), .B(n4745), .Y(n391) );
  INVX1 U3300 ( .A(n391), .Y(n3439) );
  AND2X1 U3301 ( .A(fifo_array[211]), .B(n4745), .Y(n379) );
  INVX1 U3302 ( .A(n379), .Y(n3440) );
  AND2X1 U3303 ( .A(fifo_array[186]), .B(n4747), .Y(n352) );
  INVX1 U3304 ( .A(n352), .Y(n3441) );
  AND2X1 U3305 ( .A(fifo_array[174]), .B(n4747), .Y(n340) );
  INVX1 U3306 ( .A(n340), .Y(n3442) );
  AND2X1 U3307 ( .A(fifo_array[153]), .B(n4749), .Y(n317) );
  INVX1 U3308 ( .A(n317), .Y(n3443) );
  AND2X1 U3309 ( .A(fifo_array[141]), .B(n4749), .Y(n305) );
  INVX1 U3310 ( .A(n305), .Y(n3444) );
  AND2X1 U3311 ( .A(fifo_array[116]), .B(n4751), .Y(n278) );
  INVX1 U3312 ( .A(n278), .Y(n3445) );
  AND2X1 U3313 ( .A(fifo_array[104]), .B(n4751), .Y(n266) );
  INVX1 U3314 ( .A(n266), .Y(n3446) );
  AND2X1 U3315 ( .A(fifo_array[83]), .B(n4753), .Y(n243) );
  INVX1 U3316 ( .A(n243), .Y(n3447) );
  AND2X1 U3317 ( .A(fifo_array[71]), .B(n4753), .Y(n231) );
  INVX1 U3318 ( .A(n231), .Y(n3448) );
  AND2X1 U3319 ( .A(fifo_array[43]), .B(n4755), .Y(n201) );
  INVX1 U3320 ( .A(n201), .Y(n3449) );
  AND2X1 U3321 ( .A(fifo_array[34]), .B(n4755), .Y(n192) );
  INVX1 U3322 ( .A(n192), .Y(n3450) );
  AND2X1 U3323 ( .A(fifo_array[13]), .B(n4757), .Y(n168) );
  INVX1 U3324 ( .A(n168), .Y(n3451) );
  AND2X1 U3325 ( .A(fifo_array[1]), .B(n4757), .Y(n156) );
  INVX1 U3326 ( .A(n156), .Y(n3452) );
  AND2X1 U3327 ( .A(fillcount[2]), .B(fillcount[3]), .Y(n1362) );
  INVX1 U3328 ( .A(n1362), .Y(n3453) );
  AND2X1 U3329 ( .A(put), .B(n4805), .Y(n1359) );
  INVX1 U3330 ( .A(n1359), .Y(n3454) );
  AND2X1 U3331 ( .A(n4759), .B(n4764), .Y(n4760) );
  INVX1 U3332 ( .A(n4760), .Y(n3455) );
  AND2X1 U3333 ( .A(n4758), .B(n3523), .Y(n1348) );
  INVX1 U3334 ( .A(n1348), .Y(n3456) );
  INVX1 U3335 ( .A(n1288), .Y(n3457) );
  AND2X1 U3336 ( .A(fifo_array[1071]), .B(n4695), .Y(n1269) );
  INVX1 U3337 ( .A(n1269), .Y(n3458) );
  AND2X1 U3338 ( .A(fifo_array[1059]), .B(n4695), .Y(n1257) );
  INVX1 U3339 ( .A(n1257), .Y(n3459) );
  AND2X1 U3340 ( .A(fifo_array[1036]), .B(n4697), .Y(n1233) );
  INVX1 U3341 ( .A(n1233), .Y(n3460) );
  AND2X1 U3342 ( .A(fifo_array[1024]), .B(n4697), .Y(n1221) );
  INVX1 U3343 ( .A(n1221), .Y(n3461) );
  AND2X1 U3344 ( .A(fifo_array[1001]), .B(n4699), .Y(n1197) );
  INVX1 U3345 ( .A(n1197), .Y(n3462) );
  AND2X1 U3346 ( .A(fifo_array[989]), .B(n4699), .Y(n1185) );
  INVX1 U3347 ( .A(n1185), .Y(n3463) );
  AND2X1 U3348 ( .A(fifo_array[966]), .B(n4701), .Y(n1161) );
  INVX1 U3349 ( .A(n1161), .Y(n3464) );
  AND2X1 U3350 ( .A(fifo_array[954]), .B(n4701), .Y(n1149) );
  INVX1 U3351 ( .A(n1149), .Y(n3465) );
  AND2X1 U3352 ( .A(fifo_array[931]), .B(n4703), .Y(n1125) );
  INVX1 U3353 ( .A(n1125), .Y(n3466) );
  AND2X1 U3354 ( .A(fifo_array[919]), .B(n4703), .Y(n1113) );
  INVX1 U3355 ( .A(n1113), .Y(n3467) );
  AND2X1 U3356 ( .A(fifo_array[893]), .B(n4705), .Y(n1086) );
  INVX1 U3357 ( .A(n1086), .Y(n3468) );
  AND2X1 U3358 ( .A(fifo_array[884]), .B(n4705), .Y(n1077) );
  INVX1 U3359 ( .A(n1077), .Y(n3469) );
  AND2X1 U3360 ( .A(fifo_array[873]), .B(n4707), .Y(n1065) );
  INVX1 U3361 ( .A(n1065), .Y(n3470) );
  AND2X1 U3362 ( .A(fifo_array[845]), .B(n4709), .Y(n1035) );
  INVX1 U3363 ( .A(n1035), .Y(n3471) );
  AND2X1 U3364 ( .A(fifo_array[828]), .B(n4709), .Y(n1018) );
  INVX1 U3365 ( .A(n1018), .Y(n3472) );
  AND2X1 U3366 ( .A(fifo_array[804]), .B(n4710), .Y(n993) );
  INVX1 U3367 ( .A(n993), .Y(n3473) );
  AND2X1 U3368 ( .A(fifo_array[793]), .B(n4711), .Y(n982) );
  INVX1 U3369 ( .A(n982), .Y(n3474) );
  AND2X1 U3370 ( .A(fifo_array[769]), .B(n4712), .Y(n957) );
  INVX1 U3371 ( .A(n957), .Y(n3475) );
  AND2X1 U3372 ( .A(fifo_array[758]), .B(n4713), .Y(n946) );
  INVX1 U3373 ( .A(n946), .Y(n3476) );
  AND2X1 U3374 ( .A(fifo_array[734]), .B(n4714), .Y(n921) );
  INVX1 U3375 ( .A(n921), .Y(n3477) );
  AND2X1 U3376 ( .A(fifo_array[722]), .B(n4714), .Y(n909) );
  INVX1 U3377 ( .A(n909), .Y(n3478) );
  AND2X1 U3378 ( .A(fifo_array[699]), .B(n4717), .Y(n885) );
  INVX1 U3379 ( .A(n885), .Y(n3479) );
  AND2X1 U3380 ( .A(fifo_array[687]), .B(n4716), .Y(n873) );
  INVX1 U3381 ( .A(n873), .Y(n3480) );
  AND2X1 U3382 ( .A(fifo_array[664]), .B(n4719), .Y(n849) );
  INVX1 U3383 ( .A(n849), .Y(n3481) );
  AND2X1 U3384 ( .A(fifo_array[652]), .B(n4718), .Y(n837) );
  INVX1 U3385 ( .A(n837), .Y(n3482) );
  AND2X1 U3386 ( .A(fifo_array[629]), .B(n4721), .Y(n813) );
  INVX1 U3387 ( .A(n813), .Y(n3483) );
  AND2X1 U3388 ( .A(fifo_array[617]), .B(n4720), .Y(n801) );
  INVX1 U3389 ( .A(n801), .Y(n3484) );
  AND2X1 U3390 ( .A(fifo_array[594]), .B(n4723), .Y(n777) );
  INVX1 U3391 ( .A(n777), .Y(n3485) );
  AND2X1 U3392 ( .A(fifo_array[582]), .B(n4722), .Y(n765) );
  INVX1 U3393 ( .A(n765), .Y(n3486) );
  AND2X1 U3394 ( .A(fifo_array[559]), .B(n4725), .Y(n740) );
  INVX1 U3395 ( .A(n740), .Y(n3487) );
  AND2X1 U3396 ( .A(fifo_array[547]), .B(n4724), .Y(n728) );
  INVX1 U3397 ( .A(n728), .Y(n3488) );
  AND2X1 U3398 ( .A(fifo_array[524]), .B(n4727), .Y(n704) );
  INVX1 U3399 ( .A(n704), .Y(n3489) );
  AND2X1 U3400 ( .A(fifo_array[512]), .B(n4726), .Y(n692) );
  INVX1 U3401 ( .A(n692), .Y(n3490) );
  AND2X1 U3402 ( .A(fifo_array[489]), .B(n4729), .Y(n668) );
  INVX1 U3403 ( .A(n668), .Y(n3491) );
  AND2X1 U3404 ( .A(fifo_array[477]), .B(n4728), .Y(n656) );
  INVX1 U3405 ( .A(n656), .Y(n3492) );
  AND2X1 U3406 ( .A(fifo_array[451]), .B(n4731), .Y(n629) );
  INVX1 U3407 ( .A(n629), .Y(n3493) );
  AND2X1 U3408 ( .A(fifo_array[442]), .B(n4730), .Y(n620) );
  INVX1 U3409 ( .A(n620), .Y(n3494) );
  AND2X1 U3410 ( .A(fifo_array[431]), .B(n4733), .Y(n608) );
  INVX1 U3411 ( .A(n608), .Y(n3495) );
  AND2X1 U3412 ( .A(fifo_array[403]), .B(n4734), .Y(n579) );
  INVX1 U3413 ( .A(n579), .Y(n3496) );
  AND2X1 U3414 ( .A(fifo_array[386]), .B(n4735), .Y(n562) );
  INVX1 U3415 ( .A(n562), .Y(n3497) );
  AND2X1 U3416 ( .A(fifo_array[362]), .B(n4736), .Y(n537) );
  INVX1 U3417 ( .A(n537), .Y(n3498) );
  AND2X1 U3418 ( .A(fifo_array[351]), .B(n4737), .Y(n526) );
  INVX1 U3419 ( .A(n526), .Y(n3499) );
  AND2X1 U3420 ( .A(fifo_array[327]), .B(n4738), .Y(n501) );
  INVX1 U3421 ( .A(n501), .Y(n3500) );
  AND2X1 U3422 ( .A(fifo_array[316]), .B(n4739), .Y(n490) );
  INVX1 U3423 ( .A(n490), .Y(n3501) );
  AND2X1 U3424 ( .A(fifo_array[292]), .B(n4740), .Y(n464) );
  INVX1 U3425 ( .A(n464), .Y(n3502) );
  AND2X1 U3426 ( .A(fifo_array[280]), .B(n4740), .Y(n452) );
  INVX1 U3427 ( .A(n452), .Y(n3503) );
  AND2X1 U3428 ( .A(fifo_array[257]), .B(n4743), .Y(n427) );
  INVX1 U3429 ( .A(n427), .Y(n3504) );
  AND2X1 U3430 ( .A(fifo_array[245]), .B(n4743), .Y(n415) );
  INVX1 U3431 ( .A(n415), .Y(n3505) );
  AND2X1 U3432 ( .A(fifo_array[222]), .B(n4745), .Y(n390) );
  INVX1 U3433 ( .A(n390), .Y(n3506) );
  AND2X1 U3434 ( .A(fifo_array[210]), .B(n4745), .Y(n378) );
  INVX1 U3435 ( .A(n378), .Y(n3507) );
  AND2X1 U3436 ( .A(fifo_array[187]), .B(n4747), .Y(n353) );
  INVX1 U3437 ( .A(n353), .Y(n3508) );
  AND2X1 U3438 ( .A(fifo_array[175]), .B(n4747), .Y(n341) );
  INVX1 U3439 ( .A(n341), .Y(n3509) );
  AND2X1 U3440 ( .A(fifo_array[152]), .B(n4749), .Y(n316) );
  INVX1 U3441 ( .A(n316), .Y(n3510) );
  AND2X1 U3442 ( .A(fifo_array[140]), .B(n4749), .Y(n304) );
  INVX1 U3443 ( .A(n304), .Y(n3511) );
  AND2X1 U3444 ( .A(fifo_array[117]), .B(n4751), .Y(n279) );
  INVX1 U3445 ( .A(n279), .Y(n3512) );
  AND2X1 U3446 ( .A(fifo_array[105]), .B(n4751), .Y(n267) );
  INVX1 U3447 ( .A(n267), .Y(n3513) );
  AND2X1 U3448 ( .A(fifo_array[82]), .B(n4753), .Y(n242) );
  INVX1 U3449 ( .A(n242), .Y(n3514) );
  AND2X1 U3450 ( .A(fifo_array[70]), .B(n4753), .Y(n230) );
  INVX1 U3451 ( .A(n230), .Y(n3515) );
  AND2X1 U3452 ( .A(fifo_array[47]), .B(n4755), .Y(n205) );
  INVX1 U3453 ( .A(n205), .Y(n3516) );
  AND2X1 U3454 ( .A(fifo_array[35]), .B(n4755), .Y(n193) );
  INVX1 U3455 ( .A(n193), .Y(n3517) );
  AND2X1 U3456 ( .A(fifo_array[9]), .B(n4757), .Y(n164) );
  INVX1 U3457 ( .A(n164), .Y(n3518) );
  AND2X1 U3458 ( .A(fifo_array[0]), .B(n4757), .Y(n155) );
  INVX1 U3459 ( .A(n155), .Y(n3519) );
  AND2X1 U3460 ( .A(n4813), .B(n4806), .Y(n1352) );
  INVX1 U3461 ( .A(n1352), .Y(n3520) );
  AND2X1 U3462 ( .A(n4814), .B(n95), .Y(n4759) );
  INVX1 U3463 ( .A(n4759), .Y(n3521) );
  AND2X1 U3464 ( .A(n4760), .B(n4763), .Y(n4761) );
  INVX1 U3465 ( .A(n4761), .Y(n3522) );
  BUFX2 U3466 ( .A(n1344), .Y(n3523) );
  AND2X1 U3467 ( .A(n1288), .B(n4758), .Y(n1286) );
  INVX1 U3468 ( .A(n1286), .Y(n3524) );
  INVX1 U3469 ( .A(n4583), .Y(n4632) );
  INVX1 U3470 ( .A(n4586), .Y(n4631) );
  INVX1 U3471 ( .A(n4584), .Y(n4630) );
  INVX1 U3472 ( .A(n4582), .Y(n4629) );
  INVX1 U3473 ( .A(n4580), .Y(n4628) );
  INVX1 U3474 ( .A(n4581), .Y(n4627) );
  INVX1 U3475 ( .A(n4580), .Y(n4626) );
  INVX1 U3476 ( .A(n4580), .Y(n4625) );
  INVX1 U3477 ( .A(n4580), .Y(n4624) );
  INVX1 U3478 ( .A(n4581), .Y(n4623) );
  INVX1 U3479 ( .A(n4581), .Y(n4622) );
  INVX1 U3480 ( .A(n4581), .Y(n4621) );
  INVX1 U3481 ( .A(n4582), .Y(n4620) );
  INVX1 U3482 ( .A(n4582), .Y(n4619) );
  INVX1 U3483 ( .A(n4582), .Y(n4618) );
  INVX1 U3484 ( .A(n4581), .Y(n4617) );
  INVX1 U3485 ( .A(n4580), .Y(n4616) );
  INVX1 U3486 ( .A(n4582), .Y(n4615) );
  INVX1 U3487 ( .A(n4586), .Y(n4614) );
  INVX1 U3488 ( .A(n4584), .Y(n4613) );
  INVX1 U3489 ( .A(n4580), .Y(n4612) );
  INVX1 U3490 ( .A(n4581), .Y(n4611) );
  INVX1 U3491 ( .A(n4580), .Y(n4610) );
  INVX1 U3492 ( .A(n4582), .Y(n4609) );
  INVX1 U3493 ( .A(n4583), .Y(n4608) );
  INVX1 U3494 ( .A(n4583), .Y(n4607) );
  INVX1 U3495 ( .A(n4583), .Y(n4606) );
  INVX1 U3496 ( .A(n4584), .Y(n4605) );
  INVX1 U3497 ( .A(n4584), .Y(n4604) );
  INVX1 U3498 ( .A(n4584), .Y(n4603) );
  INVX1 U3499 ( .A(n4585), .Y(n4602) );
  INVX1 U3500 ( .A(n4585), .Y(n4601) );
  INVX1 U3501 ( .A(n4585), .Y(n4600) );
  INVX1 U3502 ( .A(n4586), .Y(n4599) );
  INVX1 U3503 ( .A(n4586), .Y(n4598) );
  INVX1 U3504 ( .A(n4586), .Y(n4597) );
  INVX1 U3505 ( .A(n4587), .Y(n4596) );
  INVX1 U3506 ( .A(n4587), .Y(n4595) );
  INVX1 U3507 ( .A(n4587), .Y(n4594) );
  INVX1 U3508 ( .A(n4588), .Y(n4593) );
  INVX1 U3509 ( .A(n4588), .Y(n4592) );
  INVX1 U3510 ( .A(n4588), .Y(n4591) );
  INVX1 U3511 ( .A(n4587), .Y(n4590) );
  INVX1 U3512 ( .A(n4588), .Y(n4589) );
  INVX1 U3513 ( .A(n3525), .Y(n4691) );
  INVX1 U3514 ( .A(n1251), .Y(n4695) );
  INVX1 U3515 ( .A(n1251), .Y(n4694) );
  INVX1 U3516 ( .A(n19), .Y(n4580) );
  INVX1 U3517 ( .A(n19), .Y(n4581) );
  INVX1 U3518 ( .A(n19), .Y(n4582) );
  INVX1 U3519 ( .A(n4634), .Y(n4583) );
  INVX1 U3520 ( .A(n4634), .Y(n4584) );
  INVX1 U3521 ( .A(n4634), .Y(n4585) );
  INVX1 U3522 ( .A(n4634), .Y(n4586) );
  INVX1 U3523 ( .A(n19), .Y(n4587) );
  INVX1 U3524 ( .A(n19), .Y(n4588) );
  AND2X1 U3525 ( .A(n1354), .B(n1295), .Y(n1298) );
  AND2X1 U3526 ( .A(n1355), .B(n1295), .Y(n1297) );
  AND2X1 U3527 ( .A(n3525), .B(n4758), .Y(n1305) );
  INVX1 U3528 ( .A(n4693), .Y(n4692) );
  INVX1 U3529 ( .A(n549), .Y(n4735) );
  INVX1 U3530 ( .A(n619), .Y(n4731) );
  INVX1 U3531 ( .A(n654), .Y(n4729) );
  INVX1 U3532 ( .A(n689), .Y(n4727) );
  INVX1 U3533 ( .A(n830), .Y(n4719) );
  INVX1 U3534 ( .A(n900), .Y(n4715) );
  INVX1 U3535 ( .A(n935), .Y(n4713) );
  INVX1 U3536 ( .A(n970), .Y(n4711) );
  INVX1 U3537 ( .A(n1111), .Y(n4703) );
  INVX1 U3538 ( .A(n1181), .Y(n4699) );
  INVX1 U3539 ( .A(n1216), .Y(n4697) );
  INVX1 U3540 ( .A(n443), .Y(n4741) );
  INVX1 U3541 ( .A(n479), .Y(n4739) );
  INVX1 U3542 ( .A(n724), .Y(n4725) );
  INVX1 U3543 ( .A(n760), .Y(n4723) );
  INVX1 U3544 ( .A(n1005), .Y(n4709) );
  INVX1 U3545 ( .A(n1041), .Y(n4707) );
  INVX1 U3546 ( .A(n514), .Y(n4737) );
  INVX1 U3547 ( .A(n584), .Y(n4733) );
  INVX1 U3548 ( .A(n795), .Y(n4721) );
  INVX1 U3549 ( .A(n865), .Y(n4717) );
  INVX1 U3550 ( .A(n1076), .Y(n4705) );
  INVX1 U3551 ( .A(n1146), .Y(n4701) );
  INVX1 U3552 ( .A(n549), .Y(n4734) );
  INVX1 U3553 ( .A(n619), .Y(n4730) );
  INVX1 U3554 ( .A(n654), .Y(n4728) );
  INVX1 U3555 ( .A(n689), .Y(n4726) );
  INVX1 U3556 ( .A(n830), .Y(n4718) );
  INVX1 U3557 ( .A(n900), .Y(n4714) );
  INVX1 U3558 ( .A(n935), .Y(n4712) );
  INVX1 U3559 ( .A(n970), .Y(n4710) );
  INVX1 U3560 ( .A(n1111), .Y(n4702) );
  INVX1 U3561 ( .A(n1181), .Y(n4698) );
  INVX1 U3562 ( .A(n1216), .Y(n4696) );
  INVX1 U3563 ( .A(n443), .Y(n4740) );
  INVX1 U3564 ( .A(n479), .Y(n4738) );
  INVX1 U3565 ( .A(n724), .Y(n4724) );
  INVX1 U3566 ( .A(n760), .Y(n4722) );
  INVX1 U3567 ( .A(n1005), .Y(n4708) );
  INVX1 U3568 ( .A(n1041), .Y(n4706) );
  INVX1 U3569 ( .A(n514), .Y(n4736) );
  INVX1 U3570 ( .A(n584), .Y(n4732) );
  INVX1 U3571 ( .A(n795), .Y(n4720) );
  INVX1 U3572 ( .A(n865), .Y(n4716) );
  INVX1 U3573 ( .A(n1076), .Y(n4704) );
  INVX1 U3574 ( .A(n1146), .Y(n4700) );
  INVX1 U3575 ( .A(n154), .Y(n4757) );
  INVX1 U3576 ( .A(n191), .Y(n4755) );
  INVX1 U3577 ( .A(n227), .Y(n4753) );
  INVX1 U3578 ( .A(n263), .Y(n4751) );
  INVX1 U3579 ( .A(n299), .Y(n4749) );
  INVX1 U3580 ( .A(n335), .Y(n4747) );
  INVX1 U3581 ( .A(n371), .Y(n4745) );
  INVX1 U3582 ( .A(n407), .Y(n4743) );
  AND2X1 U3583 ( .A(n1359), .B(n4758), .Y(n1354) );
  INVX1 U3584 ( .A(n191), .Y(n4754) );
  INVX1 U3585 ( .A(n227), .Y(n4752) );
  INVX1 U3586 ( .A(n263), .Y(n4750) );
  INVX1 U3587 ( .A(n299), .Y(n4748) );
  INVX1 U3588 ( .A(n335), .Y(n4746) );
  INVX1 U3589 ( .A(n371), .Y(n4744) );
  INVX1 U3590 ( .A(n407), .Y(n4742) );
  INVX1 U3591 ( .A(n154), .Y(n4756) );
  INVX1 U3592 ( .A(n4653), .Y(n4651) );
  INVX1 U3593 ( .A(n4653), .Y(n4650) );
  INVX1 U3594 ( .A(n4653), .Y(n4649) );
  INVX1 U3595 ( .A(n4653), .Y(n4648) );
  INVX1 U3596 ( .A(n4653), .Y(n4647) );
  INVX1 U3597 ( .A(n4653), .Y(n4646) );
  INVX1 U3598 ( .A(n4653), .Y(n4645) );
  INVX1 U3599 ( .A(n4653), .Y(n4644) );
  INVX1 U3600 ( .A(n4653), .Y(n4643) );
  INVX1 U3601 ( .A(n4653), .Y(n4642) );
  INVX1 U3602 ( .A(n4653), .Y(n4641) );
  INVX1 U3603 ( .A(n4653), .Y(n4640) );
  INVX1 U3604 ( .A(n4653), .Y(n4639) );
  INVX1 U3605 ( .A(n4653), .Y(n4638) );
  INVX1 U3606 ( .A(n4653), .Y(n4637) );
  INVX1 U3607 ( .A(n4653), .Y(n4636) );
  INVX1 U3608 ( .A(n4653), .Y(n4635) );
  INVX1 U3609 ( .A(n4656), .Y(n4655) );
  INVX1 U3610 ( .A(n4656), .Y(n4654) );
  INVX1 U3611 ( .A(n4653), .Y(n4652) );
  INVX1 U3612 ( .A(n4587), .Y(n4633) );
  INVX1 U3613 ( .A(n4588), .Y(n4634) );
  INVX1 U3614 ( .A(n3525), .Y(n4693) );
  INVX1 U3615 ( .A(reset), .Y(n4758) );
  INVX1 U3616 ( .A(n82), .Y(n4800) );
  INVX1 U3617 ( .A(n3523), .Y(n4765) );
  INVX1 U3618 ( .A(data_in[0]), .Y(n4664) );
  INVX1 U3619 ( .A(data_in[1]), .Y(n4663) );
  INVX1 U3620 ( .A(data_in[2]), .Y(n4662) );
  INVX1 U3621 ( .A(data_in[3]), .Y(n4661) );
  INVX1 U3622 ( .A(data_in[4]), .Y(n4660) );
  INVX1 U3623 ( .A(data_in[5]), .Y(n4690) );
  INVX1 U3624 ( .A(data_in[6]), .Y(n4689) );
  INVX1 U3625 ( .A(data_in[7]), .Y(n4688) );
  INVX1 U3626 ( .A(data_in[8]), .Y(n4687) );
  INVX1 U3627 ( .A(data_in[9]), .Y(n4686) );
  INVX1 U3628 ( .A(data_in[10]), .Y(n4685) );
  INVX1 U3629 ( .A(data_in[11]), .Y(n4684) );
  INVX1 U3630 ( .A(data_in[12]), .Y(n4683) );
  INVX1 U3631 ( .A(data_in[13]), .Y(n4682) );
  INVX1 U3632 ( .A(data_in[14]), .Y(n4681) );
  INVX1 U3633 ( .A(data_in[15]), .Y(n4680) );
  INVX1 U3634 ( .A(data_in[16]), .Y(n4679) );
  INVX1 U3635 ( .A(data_in[17]), .Y(n4678) );
  INVX1 U3636 ( .A(data_in[18]), .Y(n4677) );
  INVX1 U3637 ( .A(data_in[19]), .Y(n4676) );
  INVX1 U3638 ( .A(data_in[20]), .Y(n4675) );
  INVX1 U3639 ( .A(data_in[21]), .Y(n4674) );
  INVX1 U3640 ( .A(data_in[22]), .Y(n4673) );
  INVX1 U3641 ( .A(data_in[23]), .Y(n4672) );
  INVX1 U3642 ( .A(data_in[24]), .Y(n4671) );
  INVX1 U3643 ( .A(data_in[25]), .Y(n4670) );
  INVX1 U3644 ( .A(data_in[26]), .Y(n4669) );
  INVX1 U3645 ( .A(data_in[27]), .Y(n4668) );
  INVX1 U3646 ( .A(data_in[28]), .Y(n4667) );
  INVX1 U3647 ( .A(data_in[29]), .Y(n4666) );
  INVX1 U3648 ( .A(data_in[30]), .Y(n4665) );
  INVX1 U3649 ( .A(data_in[31]), .Y(n4659) );
  INVX1 U3650 ( .A(data_in[32]), .Y(n4658) );
  INVX1 U3651 ( .A(data_in[33]), .Y(n4657) );
  INVX1 U3652 ( .A(n91), .Y(n4804) );
  INVX1 U3653 ( .A(n78), .Y(n4796) );
  INVX1 U3654 ( .A(n4576), .Y(n27) );
  INVX1 U3655 ( .A(n77), .Y(n4795) );
  INVX1 U3656 ( .A(n4575), .Y(n28) );
  INVX1 U3657 ( .A(n72), .Y(n4794) );
  INVX1 U3658 ( .A(n4574), .Y(n29) );
  INVX1 U3659 ( .A(n67), .Y(n4793) );
  INVX1 U3660 ( .A(n4573), .Y(n30) );
  INVX1 U3661 ( .A(n66), .Y(n4792) );
  INVX1 U3662 ( .A(n4572), .Y(n31) );
  INVX1 U3663 ( .A(n65), .Y(n4791) );
  INVX1 U3664 ( .A(n4571), .Y(n32) );
  INVX1 U3665 ( .A(n64), .Y(n4790) );
  INVX1 U3666 ( .A(n4570), .Y(n33) );
  INVX1 U3667 ( .A(n63), .Y(n4789) );
  INVX1 U3668 ( .A(n4569), .Y(n34) );
  INVX1 U3669 ( .A(n62), .Y(n4788) );
  INVX1 U3670 ( .A(n4568), .Y(n35) );
  INVX1 U3671 ( .A(n61), .Y(n4787) );
  INVX1 U3672 ( .A(n4567), .Y(n36) );
  INVX1 U3673 ( .A(n60), .Y(n4786) );
  INVX1 U3674 ( .A(n4566), .Y(n37) );
  INVX1 U3675 ( .A(n59), .Y(n4785) );
  INVX1 U3676 ( .A(n4565), .Y(n38) );
  INVX1 U3677 ( .A(n58), .Y(n4784) );
  INVX1 U3678 ( .A(n4564), .Y(n39) );
  INVX1 U3679 ( .A(n18), .Y(n4783) );
  INVX1 U3680 ( .A(n4563), .Y(n40) );
  INVX1 U3681 ( .A(n17), .Y(n4782) );
  INVX1 U3682 ( .A(n4562), .Y(n41) );
  INVX1 U3683 ( .A(n16), .Y(n4781) );
  INVX1 U3684 ( .A(n4561), .Y(n42) );
  INVX1 U3685 ( .A(n15), .Y(n4780) );
  INVX1 U3686 ( .A(n4560), .Y(n43) );
  INVX1 U3687 ( .A(n14), .Y(n4779) );
  INVX1 U3688 ( .A(n4559), .Y(n44) );
  INVX1 U3689 ( .A(n13), .Y(n4778) );
  INVX1 U3690 ( .A(n4558), .Y(n45) );
  INVX1 U3691 ( .A(n12), .Y(n4777) );
  INVX1 U3692 ( .A(n4557), .Y(n46) );
  INVX1 U3693 ( .A(n11), .Y(n4776) );
  INVX1 U3694 ( .A(n4556), .Y(n47) );
  INVX1 U3695 ( .A(n10), .Y(n4775) );
  INVX1 U3696 ( .A(n4555), .Y(n48) );
  INVX1 U3697 ( .A(n9), .Y(n4774) );
  INVX1 U3698 ( .A(n4554), .Y(n49) );
  INVX1 U3699 ( .A(n8), .Y(n4773) );
  INVX1 U3700 ( .A(n4553), .Y(n50) );
  INVX1 U3701 ( .A(n7), .Y(n4772) );
  INVX1 U3702 ( .A(n4552), .Y(n51) );
  INVX1 U3703 ( .A(n6), .Y(n4771) );
  INVX1 U3704 ( .A(n4551), .Y(n52) );
  INVX1 U3705 ( .A(n80), .Y(n4798) );
  INVX1 U3706 ( .A(n4578), .Y(n25) );
  INVX1 U3707 ( .A(n90), .Y(n4803) );
  INVX1 U3708 ( .A(n89), .Y(n4802) );
  INVX1 U3709 ( .A(n83), .Y(n4801) );
  INVX1 U3710 ( .A(n3), .Y(n4768) );
  INVX1 U3711 ( .A(n4548), .Y(n55) );
  INVX1 U3712 ( .A(n2), .Y(n4767) );
  INVX1 U3713 ( .A(n4547), .Y(n56) );
  INVX1 U3714 ( .A(n1), .Y(n4766) );
  INVX1 U3715 ( .A(n4546), .Y(n57) );
  INVX1 U3716 ( .A(n4), .Y(n4769) );
  INVX1 U3717 ( .A(n4549), .Y(n54) );
  INVX1 U3718 ( .A(n5), .Y(n4770) );
  INVX1 U3719 ( .A(n4550), .Y(n53) );
  INVX1 U3720 ( .A(n81), .Y(n4799) );
  INVX1 U3721 ( .A(n4579), .Y(n24) );
  INVX1 U3722 ( .A(n79), .Y(n4797) );
  INVX1 U3723 ( .A(n4577), .Y(n26) );
  INVX1 U3724 ( .A(empty), .Y(n4807) );
  INVX1 U3725 ( .A(full), .Y(n4805) );
  INVX1 U3726 ( .A(wr_ptr[2]), .Y(n4810) );
  INVX1 U3727 ( .A(wr_ptr[0]), .Y(n4808) );
  INVX1 U3728 ( .A(wr_ptr[1]), .Y(n4809) );
  INVX1 U3729 ( .A(n20), .Y(n4653) );
  INVX1 U3730 ( .A(wr_ptr[4]), .Y(n4812) );
  INVX1 U3731 ( .A(wr_ptr[3]), .Y(n4811) );
  INVX1 U3732 ( .A(n21), .Y(n4656) );
  INVX1 U3733 ( .A(fillcount[4]), .Y(n4813) );
  INVX1 U3734 ( .A(fillcount[0]), .Y(n95) );
  INVX1 U3735 ( .A(fillcount[5]), .Y(n4806) );
  INVX1 U3736 ( .A(fillcount[2]), .Y(n4764) );
  INVX1 U3737 ( .A(fillcount[3]), .Y(n4763) );
  INVX1 U3738 ( .A(fillcount[1]), .Y(n4814) );
  AND2X1 U3739 ( .A(n4814), .B(fillcount[0]), .Y(n1350) );
  MUX2X1 U3740 ( .B(n3527), .A(n3528), .S(n20), .Y(n3526) );
  MUX2X1 U3741 ( .B(n3530), .A(n3531), .S(n20), .Y(n3529) );
  MUX2X1 U3742 ( .B(n3533), .A(n3534), .S(n20), .Y(n3532) );
  MUX2X1 U3743 ( .B(n3536), .A(n3537), .S(n20), .Y(n3535) );
  MUX2X1 U3744 ( .B(n3539), .A(n3540), .S(n22), .Y(n3538) );
  MUX2X1 U3745 ( .B(n3542), .A(n3543), .S(n20), .Y(n3541) );
  MUX2X1 U3746 ( .B(n3545), .A(n3546), .S(n20), .Y(n3544) );
  MUX2X1 U3747 ( .B(n3548), .A(n3549), .S(n20), .Y(n3547) );
  MUX2X1 U3748 ( .B(n3551), .A(n3552), .S(n4635), .Y(n3550) );
  MUX2X1 U3749 ( .B(n3554), .A(n3555), .S(n22), .Y(n3553) );
  MUX2X1 U3750 ( .B(n3557), .A(n3558), .S(n4635), .Y(n3556) );
  MUX2X1 U3751 ( .B(n3560), .A(n3561), .S(n4635), .Y(n3559) );
  MUX2X1 U3752 ( .B(n3563), .A(n3564), .S(n4635), .Y(n3562) );
  MUX2X1 U3753 ( .B(n3566), .A(n3567), .S(n4635), .Y(n3565) );
  MUX2X1 U3754 ( .B(n3569), .A(n3570), .S(n22), .Y(n3568) );
  MUX2X1 U3755 ( .B(n3572), .A(n3573), .S(n4635), .Y(n3571) );
  MUX2X1 U3756 ( .B(n3575), .A(n3576), .S(n4635), .Y(n3574) );
  MUX2X1 U3757 ( .B(n3578), .A(n3579), .S(n4635), .Y(n3577) );
  MUX2X1 U3758 ( .B(n3581), .A(n3582), .S(n4635), .Y(n3580) );
  MUX2X1 U3759 ( .B(n3584), .A(n3585), .S(n22), .Y(n3583) );
  MUX2X1 U3760 ( .B(n3587), .A(n3588), .S(n4635), .Y(n3586) );
  MUX2X1 U3761 ( .B(n3590), .A(n3591), .S(n4635), .Y(n3589) );
  MUX2X1 U3762 ( .B(n3593), .A(n3594), .S(n4635), .Y(n3592) );
  MUX2X1 U3763 ( .B(n3596), .A(n3597), .S(n4635), .Y(n3595) );
  MUX2X1 U3764 ( .B(n3599), .A(n3600), .S(n22), .Y(n3598) );
  MUX2X1 U3765 ( .B(n3602), .A(n3603), .S(n4636), .Y(n3601) );
  MUX2X1 U3766 ( .B(n3605), .A(n3606), .S(n4636), .Y(n3604) );
  MUX2X1 U3767 ( .B(n3608), .A(n3609), .S(n4636), .Y(n3607) );
  MUX2X1 U3768 ( .B(n3611), .A(n3612), .S(n4636), .Y(n3610) );
  MUX2X1 U3769 ( .B(n3614), .A(n3615), .S(n22), .Y(n3613) );
  MUX2X1 U3770 ( .B(n3617), .A(n3618), .S(n4636), .Y(n3616) );
  MUX2X1 U3771 ( .B(n3620), .A(n3621), .S(n4636), .Y(n3619) );
  MUX2X1 U3772 ( .B(n3623), .A(n3624), .S(n4636), .Y(n3622) );
  MUX2X1 U3773 ( .B(n3626), .A(n3627), .S(n4636), .Y(n3625) );
  MUX2X1 U3774 ( .B(n3629), .A(n3630), .S(n22), .Y(n3628) );
  MUX2X1 U3775 ( .B(n3632), .A(n3633), .S(n4636), .Y(n3631) );
  MUX2X1 U3776 ( .B(n3635), .A(n3636), .S(n4636), .Y(n3634) );
  MUX2X1 U3777 ( .B(n3638), .A(n3639), .S(n4636), .Y(n3637) );
  MUX2X1 U3778 ( .B(n3641), .A(n3642), .S(n4636), .Y(n3640) );
  MUX2X1 U3779 ( .B(n3644), .A(n3645), .S(n22), .Y(n3643) );
  MUX2X1 U3780 ( .B(n3647), .A(n3648), .S(n4637), .Y(n3646) );
  MUX2X1 U3781 ( .B(n3650), .A(n3651), .S(n4637), .Y(n3649) );
  MUX2X1 U3782 ( .B(n3653), .A(n3654), .S(n4637), .Y(n3652) );
  MUX2X1 U3783 ( .B(n3656), .A(n3657), .S(n4637), .Y(n3655) );
  MUX2X1 U3784 ( .B(n3659), .A(n3660), .S(n22), .Y(n3658) );
  MUX2X1 U3785 ( .B(n3662), .A(n3663), .S(n4637), .Y(n3661) );
  MUX2X1 U3786 ( .B(n3665), .A(n3666), .S(n4637), .Y(n3664) );
  MUX2X1 U3787 ( .B(n3668), .A(n3669), .S(n4637), .Y(n3667) );
  MUX2X1 U3788 ( .B(n3671), .A(n3672), .S(n4637), .Y(n3670) );
  MUX2X1 U3789 ( .B(n3674), .A(n3675), .S(n22), .Y(n3673) );
  MUX2X1 U3790 ( .B(n3677), .A(n3678), .S(n4637), .Y(n3676) );
  MUX2X1 U3791 ( .B(n3680), .A(n3681), .S(n4637), .Y(n3679) );
  MUX2X1 U3792 ( .B(n3683), .A(n3684), .S(n4637), .Y(n3682) );
  MUX2X1 U3793 ( .B(n3686), .A(n3687), .S(n4637), .Y(n3685) );
  MUX2X1 U3794 ( .B(n3689), .A(n3690), .S(n22), .Y(n3688) );
  MUX2X1 U3795 ( .B(n3692), .A(n3693), .S(n4638), .Y(n3691) );
  MUX2X1 U3796 ( .B(n3695), .A(n3696), .S(n4638), .Y(n3694) );
  MUX2X1 U3797 ( .B(n3698), .A(n3699), .S(n4638), .Y(n3697) );
  MUX2X1 U3798 ( .B(n3701), .A(n3702), .S(n4638), .Y(n3700) );
  MUX2X1 U3799 ( .B(n3704), .A(n3705), .S(n22), .Y(n3703) );
  MUX2X1 U3800 ( .B(n3707), .A(n3708), .S(n4638), .Y(n3706) );
  MUX2X1 U3801 ( .B(n3710), .A(n3711), .S(n4638), .Y(n3709) );
  MUX2X1 U3802 ( .B(n3713), .A(n3714), .S(n4638), .Y(n3712) );
  MUX2X1 U3803 ( .B(n3716), .A(n3717), .S(n4638), .Y(n3715) );
  MUX2X1 U3804 ( .B(n3719), .A(n3720), .S(n22), .Y(n3718) );
  MUX2X1 U3805 ( .B(n3722), .A(n3723), .S(n4638), .Y(n3721) );
  MUX2X1 U3806 ( .B(n3725), .A(n3726), .S(n4638), .Y(n3724) );
  MUX2X1 U3807 ( .B(n3728), .A(n3729), .S(n4638), .Y(n3727) );
  MUX2X1 U3808 ( .B(n3731), .A(n3732), .S(n4638), .Y(n3730) );
  MUX2X1 U3809 ( .B(n3734), .A(n3735), .S(n22), .Y(n3733) );
  MUX2X1 U3810 ( .B(n3737), .A(n3738), .S(n4639), .Y(n3736) );
  MUX2X1 U3811 ( .B(n3740), .A(n3741), .S(n4639), .Y(n3739) );
  MUX2X1 U3812 ( .B(n3743), .A(n3744), .S(n4639), .Y(n3742) );
  MUX2X1 U3813 ( .B(n3746), .A(n3747), .S(n4639), .Y(n3745) );
  MUX2X1 U3814 ( .B(n3749), .A(n3750), .S(n22), .Y(n3748) );
  MUX2X1 U3815 ( .B(n3752), .A(n3753), .S(n4639), .Y(n3751) );
  MUX2X1 U3816 ( .B(n3755), .A(n3756), .S(n4639), .Y(n3754) );
  MUX2X1 U3817 ( .B(n3758), .A(n3759), .S(n4639), .Y(n3757) );
  MUX2X1 U3818 ( .B(n3761), .A(n3762), .S(n4639), .Y(n3760) );
  MUX2X1 U3819 ( .B(n3764), .A(n3765), .S(n22), .Y(n3763) );
  MUX2X1 U3820 ( .B(n3767), .A(n3768), .S(n4639), .Y(n3766) );
  MUX2X1 U3821 ( .B(n3770), .A(n3771), .S(n4639), .Y(n3769) );
  MUX2X1 U3822 ( .B(n3773), .A(n3774), .S(n4639), .Y(n3772) );
  MUX2X1 U3823 ( .B(n3776), .A(n3777), .S(n4639), .Y(n3775) );
  MUX2X1 U3824 ( .B(n3779), .A(n3780), .S(n22), .Y(n3778) );
  MUX2X1 U3825 ( .B(n3782), .A(n3783), .S(n4640), .Y(n3781) );
  MUX2X1 U3826 ( .B(n3785), .A(n3786), .S(n4640), .Y(n3784) );
  MUX2X1 U3827 ( .B(n3788), .A(n3789), .S(n4640), .Y(n3787) );
  MUX2X1 U3828 ( .B(n3791), .A(n3792), .S(n4640), .Y(n3790) );
  MUX2X1 U3829 ( .B(n3794), .A(n3795), .S(n22), .Y(n3793) );
  MUX2X1 U3830 ( .B(n3797), .A(n3798), .S(n4640), .Y(n3796) );
  MUX2X1 U3831 ( .B(n3800), .A(n3801), .S(n4640), .Y(n3799) );
  MUX2X1 U3832 ( .B(n3803), .A(n3804), .S(n4640), .Y(n3802) );
  MUX2X1 U3833 ( .B(n3806), .A(n3807), .S(n4640), .Y(n3805) );
  MUX2X1 U3834 ( .B(n3809), .A(n3810), .S(n22), .Y(n3808) );
  MUX2X1 U3835 ( .B(n3812), .A(n3813), .S(n4640), .Y(n3811) );
  MUX2X1 U3836 ( .B(n3815), .A(n3816), .S(n4640), .Y(n3814) );
  MUX2X1 U3837 ( .B(n3818), .A(n3819), .S(n4640), .Y(n3817) );
  MUX2X1 U3838 ( .B(n3821), .A(n3822), .S(n4640), .Y(n3820) );
  MUX2X1 U3839 ( .B(n3824), .A(n3825), .S(n22), .Y(n3823) );
  MUX2X1 U3840 ( .B(n3827), .A(n3828), .S(n4641), .Y(n3826) );
  MUX2X1 U3841 ( .B(n3830), .A(n3831), .S(n4641), .Y(n3829) );
  MUX2X1 U3842 ( .B(n3833), .A(n3834), .S(n4641), .Y(n3832) );
  MUX2X1 U3843 ( .B(n3836), .A(n3837), .S(n4641), .Y(n3835) );
  MUX2X1 U3844 ( .B(n3839), .A(n3840), .S(n22), .Y(n3838) );
  MUX2X1 U3845 ( .B(n3842), .A(n3843), .S(n4641), .Y(n3841) );
  MUX2X1 U3846 ( .B(n3845), .A(n3846), .S(n4641), .Y(n3844) );
  MUX2X1 U3847 ( .B(n3848), .A(n3849), .S(n4641), .Y(n3847) );
  MUX2X1 U3848 ( .B(n3851), .A(n3852), .S(n4641), .Y(n3850) );
  MUX2X1 U3849 ( .B(n3854), .A(n3855), .S(n22), .Y(n3853) );
  MUX2X1 U3850 ( .B(n3857), .A(n3858), .S(n4641), .Y(n3856) );
  MUX2X1 U3851 ( .B(n3860), .A(n3861), .S(n4641), .Y(n3859) );
  MUX2X1 U3852 ( .B(n3863), .A(n3864), .S(n4641), .Y(n3862) );
  MUX2X1 U3853 ( .B(n3866), .A(n3867), .S(n4641), .Y(n3865) );
  MUX2X1 U3854 ( .B(n3869), .A(n3870), .S(n22), .Y(n3868) );
  MUX2X1 U3855 ( .B(n3872), .A(n3873), .S(n4642), .Y(n3871) );
  MUX2X1 U3856 ( .B(n3875), .A(n3876), .S(n4642), .Y(n3874) );
  MUX2X1 U3857 ( .B(n3878), .A(n3879), .S(n4642), .Y(n3877) );
  MUX2X1 U3858 ( .B(n3881), .A(n3882), .S(n4642), .Y(n3880) );
  MUX2X1 U3859 ( .B(n3884), .A(n3885), .S(n22), .Y(n3883) );
  MUX2X1 U3860 ( .B(n3887), .A(n3888), .S(n4642), .Y(n3886) );
  MUX2X1 U3861 ( .B(n3890), .A(n3891), .S(n4642), .Y(n3889) );
  MUX2X1 U3862 ( .B(n3893), .A(n3894), .S(n4642), .Y(n3892) );
  MUX2X1 U3863 ( .B(n3896), .A(n3897), .S(n4642), .Y(n3895) );
  MUX2X1 U3864 ( .B(n3899), .A(n3900), .S(n22), .Y(n3898) );
  MUX2X1 U3865 ( .B(n3902), .A(n3903), .S(n4642), .Y(n3901) );
  MUX2X1 U3866 ( .B(n3905), .A(n3906), .S(n4642), .Y(n3904) );
  MUX2X1 U3867 ( .B(n3908), .A(n3909), .S(n4642), .Y(n3907) );
  MUX2X1 U3868 ( .B(n3911), .A(n3912), .S(n4642), .Y(n3910) );
  MUX2X1 U3869 ( .B(n3914), .A(n3915), .S(n22), .Y(n3913) );
  MUX2X1 U3870 ( .B(n3917), .A(n3918), .S(n4643), .Y(n3916) );
  MUX2X1 U3871 ( .B(n3920), .A(n3921), .S(n4643), .Y(n3919) );
  MUX2X1 U3872 ( .B(n3923), .A(n3924), .S(n4643), .Y(n3922) );
  MUX2X1 U3873 ( .B(n3926), .A(n3927), .S(n4643), .Y(n3925) );
  MUX2X1 U3874 ( .B(n3929), .A(n3930), .S(n22), .Y(n3928) );
  MUX2X1 U3875 ( .B(n3932), .A(n3933), .S(n4643), .Y(n3931) );
  MUX2X1 U3876 ( .B(n3935), .A(n3936), .S(n4643), .Y(n3934) );
  MUX2X1 U3877 ( .B(n3938), .A(n3939), .S(n4643), .Y(n3937) );
  MUX2X1 U3878 ( .B(n3941), .A(n3942), .S(n4643), .Y(n3940) );
  MUX2X1 U3879 ( .B(n3944), .A(n3945), .S(n22), .Y(n3943) );
  MUX2X1 U3880 ( .B(n3947), .A(n3948), .S(n4643), .Y(n3946) );
  MUX2X1 U3881 ( .B(n3950), .A(n3951), .S(n4643), .Y(n3949) );
  MUX2X1 U3882 ( .B(n3953), .A(n3954), .S(n4643), .Y(n3952) );
  MUX2X1 U3883 ( .B(n3956), .A(n3957), .S(n4643), .Y(n3955) );
  MUX2X1 U3884 ( .B(n3959), .A(n3960), .S(n22), .Y(n3958) );
  MUX2X1 U3885 ( .B(n3962), .A(n3963), .S(n4644), .Y(n3961) );
  MUX2X1 U3886 ( .B(n3965), .A(n3966), .S(n4644), .Y(n3964) );
  MUX2X1 U3887 ( .B(n3968), .A(n3969), .S(n4644), .Y(n3967) );
  MUX2X1 U3888 ( .B(n3971), .A(n3972), .S(n4644), .Y(n3970) );
  MUX2X1 U3889 ( .B(n3974), .A(n3975), .S(n22), .Y(n3973) );
  MUX2X1 U3890 ( .B(n3977), .A(n3978), .S(n4644), .Y(n3976) );
  MUX2X1 U3891 ( .B(n3980), .A(n3981), .S(n4644), .Y(n3979) );
  MUX2X1 U3892 ( .B(n3983), .A(n3984), .S(n4644), .Y(n3982) );
  MUX2X1 U3893 ( .B(n3986), .A(n3987), .S(n4644), .Y(n3985) );
  MUX2X1 U3894 ( .B(n3989), .A(n3990), .S(n22), .Y(n3988) );
  MUX2X1 U3895 ( .B(n3992), .A(n3993), .S(n4644), .Y(n3991) );
  MUX2X1 U3896 ( .B(n3995), .A(n3996), .S(n4644), .Y(n3994) );
  MUX2X1 U3897 ( .B(n3998), .A(n3999), .S(n4644), .Y(n3997) );
  MUX2X1 U3898 ( .B(n4001), .A(n4002), .S(n4644), .Y(n4000) );
  MUX2X1 U3899 ( .B(n4004), .A(n4005), .S(n22), .Y(n4003) );
  MUX2X1 U3900 ( .B(n4007), .A(n4008), .S(n4645), .Y(n4006) );
  MUX2X1 U3901 ( .B(n4010), .A(n4011), .S(n4645), .Y(n4009) );
  MUX2X1 U3902 ( .B(n4013), .A(n4014), .S(n4645), .Y(n4012) );
  MUX2X1 U3903 ( .B(n4016), .A(n4017), .S(n4645), .Y(n4015) );
  MUX2X1 U3904 ( .B(n4019), .A(n4020), .S(n22), .Y(n4018) );
  MUX2X1 U3905 ( .B(n4022), .A(n4023), .S(n4645), .Y(n4021) );
  MUX2X1 U3906 ( .B(n4025), .A(n4026), .S(n4645), .Y(n4024) );
  MUX2X1 U3907 ( .B(n4028), .A(n4029), .S(n4645), .Y(n4027) );
  MUX2X1 U3908 ( .B(n4031), .A(n4032), .S(n4645), .Y(n4030) );
  MUX2X1 U3909 ( .B(n4034), .A(n4035), .S(n22), .Y(n4033) );
  MUX2X1 U3910 ( .B(n4037), .A(n4038), .S(n4645), .Y(n4036) );
  MUX2X1 U3911 ( .B(n4040), .A(n4041), .S(n4645), .Y(n4039) );
  MUX2X1 U3912 ( .B(n4043), .A(n4044), .S(n4645), .Y(n4042) );
  MUX2X1 U3913 ( .B(n4046), .A(n4047), .S(n4645), .Y(n4045) );
  MUX2X1 U3914 ( .B(n4049), .A(n4050), .S(n22), .Y(n4048) );
  MUX2X1 U3915 ( .B(n4052), .A(n4053), .S(n4646), .Y(n4051) );
  MUX2X1 U3916 ( .B(n4055), .A(n4056), .S(n4646), .Y(n4054) );
  MUX2X1 U3917 ( .B(n4058), .A(n4059), .S(n4646), .Y(n4057) );
  MUX2X1 U3918 ( .B(n4061), .A(n4062), .S(n4646), .Y(n4060) );
  MUX2X1 U3919 ( .B(n4064), .A(n4065), .S(n22), .Y(n4063) );
  MUX2X1 U3920 ( .B(n4067), .A(n4068), .S(n4646), .Y(n4066) );
  MUX2X1 U3921 ( .B(n4070), .A(n4071), .S(n4646), .Y(n4069) );
  MUX2X1 U3922 ( .B(n4073), .A(n4074), .S(n4646), .Y(n4072) );
  MUX2X1 U3923 ( .B(n4076), .A(n4077), .S(n4646), .Y(n4075) );
  MUX2X1 U3924 ( .B(n4079), .A(n4080), .S(n22), .Y(n4078) );
  MUX2X1 U3925 ( .B(n4082), .A(n4083), .S(n4646), .Y(n4081) );
  MUX2X1 U3926 ( .B(n4085), .A(n4086), .S(n4646), .Y(n4084) );
  MUX2X1 U3927 ( .B(n4088), .A(n4089), .S(n4646), .Y(n4087) );
  MUX2X1 U3928 ( .B(n4091), .A(n4092), .S(n4646), .Y(n4090) );
  MUX2X1 U3929 ( .B(n4094), .A(n4095), .S(n22), .Y(n4093) );
  MUX2X1 U3930 ( .B(n4097), .A(n4098), .S(n4647), .Y(n4096) );
  MUX2X1 U3931 ( .B(n4100), .A(n4101), .S(n4647), .Y(n4099) );
  MUX2X1 U3932 ( .B(n4103), .A(n4104), .S(n4647), .Y(n4102) );
  MUX2X1 U3933 ( .B(n4106), .A(n4107), .S(n4647), .Y(n4105) );
  MUX2X1 U3934 ( .B(n4109), .A(n4110), .S(n22), .Y(n4108) );
  MUX2X1 U3935 ( .B(n4112), .A(n4113), .S(n4647), .Y(n4111) );
  MUX2X1 U3936 ( .B(n4115), .A(n4116), .S(n4647), .Y(n4114) );
  MUX2X1 U3937 ( .B(n4118), .A(n4119), .S(n4647), .Y(n4117) );
  MUX2X1 U3938 ( .B(n4121), .A(n4122), .S(n4647), .Y(n4120) );
  MUX2X1 U3939 ( .B(n4124), .A(n4125), .S(n22), .Y(n4123) );
  MUX2X1 U3940 ( .B(n4127), .A(n4128), .S(n4647), .Y(n4126) );
  MUX2X1 U3941 ( .B(n4130), .A(n4131), .S(n4647), .Y(n4129) );
  MUX2X1 U3942 ( .B(n4133), .A(n4134), .S(n4647), .Y(n4132) );
  MUX2X1 U3943 ( .B(n4136), .A(n4137), .S(n4647), .Y(n4135) );
  MUX2X1 U3944 ( .B(n4139), .A(n4140), .S(n22), .Y(n4138) );
  MUX2X1 U3945 ( .B(n4142), .A(n4143), .S(n4648), .Y(n4141) );
  MUX2X1 U3946 ( .B(n4145), .A(n4146), .S(n4648), .Y(n4144) );
  MUX2X1 U3947 ( .B(n4148), .A(n4149), .S(n4648), .Y(n4147) );
  MUX2X1 U3948 ( .B(n4151), .A(n4152), .S(n4648), .Y(n4150) );
  MUX2X1 U3949 ( .B(n4154), .A(n4155), .S(n22), .Y(n4153) );
  MUX2X1 U3950 ( .B(n4157), .A(n4158), .S(n4648), .Y(n4156) );
  MUX2X1 U3951 ( .B(n4160), .A(n4161), .S(n4648), .Y(n4159) );
  MUX2X1 U3952 ( .B(n4163), .A(n4164), .S(n4648), .Y(n4162) );
  MUX2X1 U3953 ( .B(n4166), .A(n4167), .S(n4648), .Y(n4165) );
  MUX2X1 U3954 ( .B(n4169), .A(n4170), .S(n22), .Y(n4168) );
  MUX2X1 U3955 ( .B(n4172), .A(n4173), .S(n4648), .Y(n4171) );
  MUX2X1 U3956 ( .B(n4175), .A(n4176), .S(n4648), .Y(n4174) );
  MUX2X1 U3957 ( .B(n4178), .A(n4179), .S(n4648), .Y(n4177) );
  MUX2X1 U3958 ( .B(n4181), .A(n4182), .S(n4648), .Y(n4180) );
  MUX2X1 U3959 ( .B(n4184), .A(n4185), .S(n22), .Y(n4183) );
  MUX2X1 U3960 ( .B(n4187), .A(n4188), .S(n4649), .Y(n4186) );
  MUX2X1 U3961 ( .B(n4190), .A(n4191), .S(n4649), .Y(n4189) );
  MUX2X1 U3962 ( .B(n4193), .A(n4194), .S(n4649), .Y(n4192) );
  MUX2X1 U3963 ( .B(n4196), .A(n4197), .S(n4649), .Y(n4195) );
  MUX2X1 U3964 ( .B(n4199), .A(n4200), .S(n22), .Y(n4198) );
  MUX2X1 U3965 ( .B(n4202), .A(n4203), .S(n4649), .Y(n4201) );
  MUX2X1 U3966 ( .B(n4205), .A(n4206), .S(n4649), .Y(n4204) );
  MUX2X1 U3967 ( .B(n4208), .A(n4209), .S(n4649), .Y(n4207) );
  MUX2X1 U3968 ( .B(n4211), .A(n4212), .S(n4649), .Y(n4210) );
  MUX2X1 U3969 ( .B(n4214), .A(n4215), .S(n22), .Y(n4213) );
  MUX2X1 U3970 ( .B(n4217), .A(n4218), .S(n4649), .Y(n4216) );
  MUX2X1 U3971 ( .B(n4220), .A(n4221), .S(n4649), .Y(n4219) );
  MUX2X1 U3972 ( .B(n4223), .A(n4224), .S(n4649), .Y(n4222) );
  MUX2X1 U3973 ( .B(n4226), .A(n4227), .S(n4649), .Y(n4225) );
  MUX2X1 U3974 ( .B(n4229), .A(n4230), .S(n22), .Y(n4228) );
  MUX2X1 U3975 ( .B(n4232), .A(n4233), .S(n4650), .Y(n4231) );
  MUX2X1 U3976 ( .B(n4235), .A(n4236), .S(n4650), .Y(n4234) );
  MUX2X1 U3977 ( .B(n4238), .A(n4239), .S(n4650), .Y(n4237) );
  MUX2X1 U3978 ( .B(n4241), .A(n4242), .S(n4650), .Y(n4240) );
  MUX2X1 U3979 ( .B(n4244), .A(n4245), .S(n22), .Y(n4243) );
  MUX2X1 U3980 ( .B(n4247), .A(n4248), .S(n4650), .Y(n4246) );
  MUX2X1 U3981 ( .B(n4250), .A(n4251), .S(n4650), .Y(n4249) );
  MUX2X1 U3982 ( .B(n4253), .A(n4254), .S(n4650), .Y(n4252) );
  MUX2X1 U3983 ( .B(n4256), .A(n4257), .S(n4650), .Y(n4255) );
  MUX2X1 U3984 ( .B(n4259), .A(n4260), .S(n22), .Y(n4258) );
  MUX2X1 U3985 ( .B(n4262), .A(n4263), .S(n4650), .Y(n4261) );
  MUX2X1 U3986 ( .B(n4265), .A(n4266), .S(n4650), .Y(n4264) );
  MUX2X1 U3987 ( .B(n4268), .A(n4269), .S(n4650), .Y(n4267) );
  MUX2X1 U3988 ( .B(n4271), .A(n4272), .S(n4650), .Y(n4270) );
  MUX2X1 U3989 ( .B(n4274), .A(n4275), .S(n22), .Y(n4273) );
  MUX2X1 U3990 ( .B(n4277), .A(n4278), .S(n4651), .Y(n4276) );
  MUX2X1 U3991 ( .B(n4280), .A(n4281), .S(n4651), .Y(n4279) );
  MUX2X1 U3992 ( .B(n4283), .A(n4284), .S(n4651), .Y(n4282) );
  MUX2X1 U3993 ( .B(n4286), .A(n4287), .S(n4651), .Y(n4285) );
  MUX2X1 U3994 ( .B(n4289), .A(n4290), .S(n22), .Y(n4288) );
  MUX2X1 U3995 ( .B(n4292), .A(n4293), .S(n4651), .Y(n4291) );
  MUX2X1 U3996 ( .B(n4295), .A(n4296), .S(n4651), .Y(n4294) );
  MUX2X1 U3997 ( .B(n4298), .A(n4299), .S(n4651), .Y(n4297) );
  MUX2X1 U3998 ( .B(n4301), .A(n4302), .S(n4651), .Y(n4300) );
  MUX2X1 U3999 ( .B(n4304), .A(n4305), .S(n22), .Y(n4303) );
  MUX2X1 U4000 ( .B(n4307), .A(n4308), .S(n4651), .Y(n4306) );
  MUX2X1 U4001 ( .B(n4310), .A(n4311), .S(n4651), .Y(n4309) );
  MUX2X1 U4002 ( .B(n4313), .A(n4314), .S(n4651), .Y(n4312) );
  MUX2X1 U4003 ( .B(n4316), .A(n4317), .S(n4651), .Y(n4315) );
  MUX2X1 U4004 ( .B(n4319), .A(n4320), .S(n22), .Y(n4318) );
  MUX2X1 U4005 ( .B(n4322), .A(n4323), .S(n4652), .Y(n4321) );
  MUX2X1 U4006 ( .B(n4325), .A(n4326), .S(n4652), .Y(n4324) );
  MUX2X1 U4007 ( .B(n4328), .A(n4329), .S(n4652), .Y(n4327) );
  MUX2X1 U4008 ( .B(n4331), .A(n4332), .S(n4652), .Y(n4330) );
  MUX2X1 U4009 ( .B(n4334), .A(n4335), .S(n22), .Y(n4333) );
  MUX2X1 U4010 ( .B(n4337), .A(n4338), .S(n4652), .Y(n4336) );
  MUX2X1 U4011 ( .B(n4340), .A(n4341), .S(n4652), .Y(n4339) );
  MUX2X1 U4012 ( .B(n4343), .A(n4344), .S(n4652), .Y(n4342) );
  MUX2X1 U4013 ( .B(n4346), .A(n4347), .S(n4652), .Y(n4345) );
  MUX2X1 U4014 ( .B(n4349), .A(n4350), .S(n22), .Y(n4348) );
  MUX2X1 U4015 ( .B(n4352), .A(n4353), .S(n4652), .Y(n4351) );
  MUX2X1 U4016 ( .B(n4355), .A(n4356), .S(n4652), .Y(n4354) );
  MUX2X1 U4017 ( .B(n4358), .A(n4359), .S(n4652), .Y(n4357) );
  MUX2X1 U4018 ( .B(n4361), .A(n4362), .S(n4652), .Y(n4360) );
  MUX2X1 U4019 ( .B(n4364), .A(n4365), .S(n22), .Y(n4363) );
  MUX2X1 U4020 ( .B(n4367), .A(n4368), .S(n4637), .Y(n4366) );
  MUX2X1 U4021 ( .B(n4370), .A(n4371), .S(n4637), .Y(n4369) );
  MUX2X1 U4022 ( .B(n4373), .A(n4374), .S(n4639), .Y(n4372) );
  MUX2X1 U4023 ( .B(n4376), .A(n4377), .S(n4651), .Y(n4375) );
  MUX2X1 U4024 ( .B(n4379), .A(n4380), .S(n22), .Y(n4378) );
  MUX2X1 U4025 ( .B(n4382), .A(n4383), .S(n4638), .Y(n4381) );
  MUX2X1 U4026 ( .B(n4385), .A(n4386), .S(n4652), .Y(n4384) );
  MUX2X1 U4027 ( .B(n4388), .A(n4389), .S(n4640), .Y(n4387) );
  MUX2X1 U4028 ( .B(n4391), .A(n4392), .S(n4641), .Y(n4390) );
  MUX2X1 U4029 ( .B(n4394), .A(n4395), .S(n22), .Y(n4393) );
  MUX2X1 U4030 ( .B(n4397), .A(n4398), .S(n4642), .Y(n4396) );
  MUX2X1 U4031 ( .B(n4400), .A(n4401), .S(n4646), .Y(n4399) );
  MUX2X1 U4032 ( .B(n4403), .A(n4404), .S(n4636), .Y(n4402) );
  MUX2X1 U4033 ( .B(n4406), .A(n4407), .S(n4643), .Y(n4405) );
  MUX2X1 U4034 ( .B(n4409), .A(n4410), .S(n22), .Y(n4408) );
  MUX2X1 U4035 ( .B(n4412), .A(n4413), .S(n4636), .Y(n4411) );
  MUX2X1 U4036 ( .B(n4415), .A(n4416), .S(n4648), .Y(n4414) );
  MUX2X1 U4037 ( .B(n4418), .A(n4419), .S(n4642), .Y(n4417) );
  MUX2X1 U4038 ( .B(n4421), .A(n4422), .S(n4647), .Y(n4420) );
  MUX2X1 U4039 ( .B(n4424), .A(n4425), .S(n22), .Y(n4423) );
  MUX2X1 U4040 ( .B(n4427), .A(n4428), .S(n4638), .Y(n4426) );
  MUX2X1 U4041 ( .B(n4430), .A(n4431), .S(n4649), .Y(n4429) );
  MUX2X1 U4042 ( .B(n4433), .A(n4434), .S(n4640), .Y(n4432) );
  MUX2X1 U4043 ( .B(n4436), .A(n4437), .S(n4644), .Y(n4435) );
  MUX2X1 U4044 ( .B(n4439), .A(n4440), .S(n22), .Y(n4438) );
  MUX2X1 U4045 ( .B(n4442), .A(n4443), .S(n4635), .Y(n4441) );
  MUX2X1 U4046 ( .B(n4445), .A(n4446), .S(n4645), .Y(n4444) );
  MUX2X1 U4047 ( .B(n4448), .A(n4449), .S(n4639), .Y(n4447) );
  MUX2X1 U4048 ( .B(n4451), .A(n4452), .S(n4650), .Y(n4450) );
  MUX2X1 U4049 ( .B(n4454), .A(n4455), .S(n22), .Y(n4453) );
  MUX2X1 U4050 ( .B(n4457), .A(n4458), .S(n20), .Y(n4456) );
  MUX2X1 U4051 ( .B(n4460), .A(n4461), .S(n20), .Y(n4459) );
  MUX2X1 U4052 ( .B(n4463), .A(n4464), .S(n20), .Y(n4462) );
  MUX2X1 U4053 ( .B(n4466), .A(n4467), .S(n20), .Y(n4465) );
  MUX2X1 U4054 ( .B(n4469), .A(n4470), .S(n22), .Y(n4468) );
  MUX2X1 U4055 ( .B(n4472), .A(n4473), .S(n20), .Y(n4471) );
  MUX2X1 U4056 ( .B(n4475), .A(n4476), .S(n20), .Y(n4474) );
  MUX2X1 U4057 ( .B(n4478), .A(n4479), .S(n20), .Y(n4477) );
  MUX2X1 U4058 ( .B(n4481), .A(n4482), .S(n20), .Y(n4480) );
  MUX2X1 U4059 ( .B(n4484), .A(n4485), .S(n22), .Y(n4483) );
  MUX2X1 U4060 ( .B(n4487), .A(n4488), .S(n20), .Y(n4486) );
  MUX2X1 U4061 ( .B(n4490), .A(n4491), .S(n20), .Y(n4489) );
  MUX2X1 U4062 ( .B(n4493), .A(n4494), .S(n20), .Y(n4492) );
  MUX2X1 U4063 ( .B(n4496), .A(n4497), .S(n20), .Y(n4495) );
  MUX2X1 U4064 ( .B(n4499), .A(n4500), .S(n22), .Y(n4498) );
  MUX2X1 U4065 ( .B(n4502), .A(n4503), .S(n4652), .Y(n4501) );
  MUX2X1 U4066 ( .B(n4505), .A(n4506), .S(n4650), .Y(n4504) );
  MUX2X1 U4067 ( .B(n4508), .A(n4509), .S(n4641), .Y(n4507) );
  MUX2X1 U4068 ( .B(n4511), .A(n4512), .S(n4644), .Y(n4510) );
  MUX2X1 U4069 ( .B(n4514), .A(n4515), .S(n22), .Y(n4513) );
  MUX2X1 U4070 ( .B(n4517), .A(n4518), .S(n4651), .Y(n4516) );
  MUX2X1 U4071 ( .B(n4520), .A(n4521), .S(n4648), .Y(n4519) );
  MUX2X1 U4072 ( .B(n4523), .A(n4524), .S(n4643), .Y(n4522) );
  MUX2X1 U4073 ( .B(n4526), .A(n4527), .S(n4647), .Y(n4525) );
  MUX2X1 U4074 ( .B(n4529), .A(n4530), .S(n22), .Y(n4528) );
  MUX2X1 U4075 ( .B(n4532), .A(n4533), .S(n4645), .Y(n4531) );
  MUX2X1 U4076 ( .B(n4535), .A(n4536), .S(n4649), .Y(n4534) );
  MUX2X1 U4077 ( .B(n4538), .A(n4539), .S(n4646), .Y(n4537) );
  MUX2X1 U4078 ( .B(n4541), .A(n4542), .S(n20), .Y(n4540) );
  MUX2X1 U4079 ( .B(n4544), .A(n4545), .S(n22), .Y(n4543) );
  MUX2X1 U4080 ( .B(fifo_array[1020]), .A(fifo_array[1054]), .S(n19), .Y(n3528) );
  MUX2X1 U4081 ( .B(fifo_array[952]), .A(fifo_array[986]), .S(n19), .Y(n3527)
         );
  MUX2X1 U4082 ( .B(fifo_array[884]), .A(fifo_array[918]), .S(n4633), .Y(n3531) );
  MUX2X1 U4083 ( .B(fifo_array[816]), .A(fifo_array[850]), .S(n4633), .Y(n3530) );
  MUX2X1 U4084 ( .B(n3529), .A(n3526), .S(n21), .Y(n3540) );
  MUX2X1 U4085 ( .B(fifo_array[748]), .A(fifo_array[782]), .S(n4589), .Y(n3534) );
  MUX2X1 U4086 ( .B(fifo_array[680]), .A(fifo_array[714]), .S(n4589), .Y(n3533) );
  MUX2X1 U4087 ( .B(fifo_array[612]), .A(fifo_array[646]), .S(n4589), .Y(n3537) );
  MUX2X1 U4088 ( .B(fifo_array[544]), .A(fifo_array[578]), .S(n4589), .Y(n3536) );
  MUX2X1 U4089 ( .B(n3535), .A(n3532), .S(n21), .Y(n3539) );
  MUX2X1 U4090 ( .B(fifo_array[476]), .A(fifo_array[510]), .S(n4589), .Y(n3543) );
  MUX2X1 U4091 ( .B(fifo_array[408]), .A(fifo_array[442]), .S(n4589), .Y(n3542) );
  MUX2X1 U4092 ( .B(fifo_array[340]), .A(fifo_array[374]), .S(n4589), .Y(n3546) );
  MUX2X1 U4093 ( .B(fifo_array[272]), .A(fifo_array[306]), .S(n4589), .Y(n3545) );
  MUX2X1 U4094 ( .B(n3544), .A(n3541), .S(n21), .Y(n3555) );
  MUX2X1 U4095 ( .B(fifo_array[204]), .A(fifo_array[238]), .S(n4589), .Y(n3549) );
  MUX2X1 U4096 ( .B(fifo_array[136]), .A(fifo_array[170]), .S(n4589), .Y(n3548) );
  MUX2X1 U4097 ( .B(fifo_array[68]), .A(fifo_array[102]), .S(n4589), .Y(n3552)
         );
  MUX2X1 U4098 ( .B(fifo_array[0]), .A(fifo_array[34]), .S(n4589), .Y(n3551)
         );
  MUX2X1 U4099 ( .B(n3550), .A(n3547), .S(n21), .Y(n3554) );
  MUX2X1 U4100 ( .B(n3553), .A(n3538), .S(n23), .Y(n4546) );
  MUX2X1 U4101 ( .B(fifo_array[1021]), .A(fifo_array[1055]), .S(n4590), .Y(
        n3558) );
  MUX2X1 U4102 ( .B(fifo_array[953]), .A(fifo_array[987]), .S(n4590), .Y(n3557) );
  MUX2X1 U4103 ( .B(fifo_array[885]), .A(fifo_array[919]), .S(n4590), .Y(n3561) );
  MUX2X1 U4104 ( .B(fifo_array[817]), .A(fifo_array[851]), .S(n4590), .Y(n3560) );
  MUX2X1 U4105 ( .B(n3559), .A(n3556), .S(n4654), .Y(n3570) );
  MUX2X1 U4106 ( .B(fifo_array[749]), .A(fifo_array[783]), .S(n4590), .Y(n3564) );
  MUX2X1 U4107 ( .B(fifo_array[681]), .A(fifo_array[715]), .S(n4590), .Y(n3563) );
  MUX2X1 U4108 ( .B(fifo_array[613]), .A(fifo_array[647]), .S(n4590), .Y(n3567) );
  MUX2X1 U4109 ( .B(fifo_array[545]), .A(fifo_array[579]), .S(n4590), .Y(n3566) );
  MUX2X1 U4110 ( .B(n3565), .A(n3562), .S(n4654), .Y(n3569) );
  MUX2X1 U4111 ( .B(fifo_array[477]), .A(fifo_array[511]), .S(n4590), .Y(n3573) );
  MUX2X1 U4112 ( .B(fifo_array[409]), .A(fifo_array[443]), .S(n4590), .Y(n3572) );
  MUX2X1 U4113 ( .B(fifo_array[341]), .A(fifo_array[375]), .S(n4590), .Y(n3576) );
  MUX2X1 U4114 ( .B(fifo_array[273]), .A(fifo_array[307]), .S(n4590), .Y(n3575) );
  MUX2X1 U4115 ( .B(n3574), .A(n3571), .S(n4654), .Y(n3585) );
  MUX2X1 U4116 ( .B(fifo_array[205]), .A(fifo_array[239]), .S(n4591), .Y(n3579) );
  MUX2X1 U4117 ( .B(fifo_array[137]), .A(fifo_array[171]), .S(n4591), .Y(n3578) );
  MUX2X1 U4118 ( .B(fifo_array[69]), .A(fifo_array[103]), .S(n4591), .Y(n3582)
         );
  MUX2X1 U4119 ( .B(fifo_array[1]), .A(fifo_array[35]), .S(n4591), .Y(n3581)
         );
  MUX2X1 U4120 ( .B(n3580), .A(n3577), .S(n4654), .Y(n3584) );
  MUX2X1 U4121 ( .B(n3583), .A(n3568), .S(n23), .Y(n4547) );
  MUX2X1 U4122 ( .B(fifo_array[1022]), .A(fifo_array[1056]), .S(n4591), .Y(
        n3588) );
  MUX2X1 U4123 ( .B(fifo_array[954]), .A(fifo_array[988]), .S(n4591), .Y(n3587) );
  MUX2X1 U4124 ( .B(fifo_array[886]), .A(fifo_array[920]), .S(n4591), .Y(n3591) );
  MUX2X1 U4125 ( .B(fifo_array[818]), .A(fifo_array[852]), .S(n4591), .Y(n3590) );
  MUX2X1 U4126 ( .B(n3589), .A(n3586), .S(n4654), .Y(n3600) );
  MUX2X1 U4127 ( .B(fifo_array[750]), .A(fifo_array[784]), .S(n4591), .Y(n3594) );
  MUX2X1 U4128 ( .B(fifo_array[682]), .A(fifo_array[716]), .S(n4591), .Y(n3593) );
  MUX2X1 U4129 ( .B(fifo_array[614]), .A(fifo_array[648]), .S(n4591), .Y(n3597) );
  MUX2X1 U4130 ( .B(fifo_array[546]), .A(fifo_array[580]), .S(n4591), .Y(n3596) );
  MUX2X1 U4131 ( .B(n3595), .A(n3592), .S(n4654), .Y(n3599) );
  MUX2X1 U4132 ( .B(fifo_array[478]), .A(fifo_array[512]), .S(n4592), .Y(n3603) );
  MUX2X1 U4133 ( .B(fifo_array[410]), .A(fifo_array[444]), .S(n4592), .Y(n3602) );
  MUX2X1 U4134 ( .B(fifo_array[342]), .A(fifo_array[376]), .S(n4592), .Y(n3606) );
  MUX2X1 U4135 ( .B(fifo_array[274]), .A(fifo_array[308]), .S(n4592), .Y(n3605) );
  MUX2X1 U4136 ( .B(n3604), .A(n3601), .S(n4654), .Y(n3615) );
  MUX2X1 U4137 ( .B(fifo_array[206]), .A(fifo_array[240]), .S(n4592), .Y(n3609) );
  MUX2X1 U4138 ( .B(fifo_array[138]), .A(fifo_array[172]), .S(n4592), .Y(n3608) );
  MUX2X1 U4139 ( .B(fifo_array[70]), .A(fifo_array[104]), .S(n4592), .Y(n3612)
         );
  MUX2X1 U4140 ( .B(fifo_array[2]), .A(fifo_array[36]), .S(n4592), .Y(n3611)
         );
  MUX2X1 U4141 ( .B(n3610), .A(n3607), .S(n4654), .Y(n3614) );
  MUX2X1 U4142 ( .B(n3613), .A(n3598), .S(n23), .Y(n4548) );
  MUX2X1 U4143 ( .B(fifo_array[1023]), .A(fifo_array[1057]), .S(n4592), .Y(
        n3618) );
  MUX2X1 U4144 ( .B(fifo_array[955]), .A(fifo_array[989]), .S(n4592), .Y(n3617) );
  MUX2X1 U4145 ( .B(fifo_array[887]), .A(fifo_array[921]), .S(n4592), .Y(n3621) );
  MUX2X1 U4146 ( .B(fifo_array[819]), .A(fifo_array[853]), .S(n4592), .Y(n3620) );
  MUX2X1 U4147 ( .B(n3619), .A(n3616), .S(n4654), .Y(n3630) );
  MUX2X1 U4148 ( .B(fifo_array[751]), .A(fifo_array[785]), .S(n4593), .Y(n3624) );
  MUX2X1 U4149 ( .B(fifo_array[683]), .A(fifo_array[717]), .S(n4593), .Y(n3623) );
  MUX2X1 U4150 ( .B(fifo_array[615]), .A(fifo_array[649]), .S(n4593), .Y(n3627) );
  MUX2X1 U4151 ( .B(fifo_array[547]), .A(fifo_array[581]), .S(n4593), .Y(n3626) );
  MUX2X1 U4152 ( .B(n3625), .A(n3622), .S(n4654), .Y(n3629) );
  MUX2X1 U4153 ( .B(fifo_array[479]), .A(fifo_array[513]), .S(n4593), .Y(n3633) );
  MUX2X1 U4154 ( .B(fifo_array[411]), .A(fifo_array[445]), .S(n4593), .Y(n3632) );
  MUX2X1 U4155 ( .B(fifo_array[343]), .A(fifo_array[377]), .S(n4593), .Y(n3636) );
  MUX2X1 U4156 ( .B(fifo_array[275]), .A(fifo_array[309]), .S(n4593), .Y(n3635) );
  MUX2X1 U4157 ( .B(n3634), .A(n3631), .S(n4654), .Y(n3645) );
  MUX2X1 U4158 ( .B(fifo_array[207]), .A(fifo_array[241]), .S(n4593), .Y(n3639) );
  MUX2X1 U4159 ( .B(fifo_array[139]), .A(fifo_array[173]), .S(n4593), .Y(n3638) );
  MUX2X1 U4160 ( .B(fifo_array[71]), .A(fifo_array[105]), .S(n4593), .Y(n3642)
         );
  MUX2X1 U4161 ( .B(fifo_array[3]), .A(fifo_array[37]), .S(n4593), .Y(n3641)
         );
  MUX2X1 U4162 ( .B(n3640), .A(n3637), .S(n4654), .Y(n3644) );
  MUX2X1 U4163 ( .B(n3643), .A(n3628), .S(n23), .Y(n4549) );
  MUX2X1 U4164 ( .B(fifo_array[1024]), .A(fifo_array[1058]), .S(n4594), .Y(
        n3648) );
  MUX2X1 U4165 ( .B(fifo_array[956]), .A(fifo_array[990]), .S(n4594), .Y(n3647) );
  MUX2X1 U4166 ( .B(fifo_array[888]), .A(fifo_array[922]), .S(n4594), .Y(n3651) );
  MUX2X1 U4167 ( .B(fifo_array[820]), .A(fifo_array[854]), .S(n4594), .Y(n3650) );
  MUX2X1 U4168 ( .B(n3649), .A(n3646), .S(n4655), .Y(n3660) );
  MUX2X1 U4169 ( .B(fifo_array[752]), .A(fifo_array[786]), .S(n4594), .Y(n3654) );
  MUX2X1 U4170 ( .B(fifo_array[684]), .A(fifo_array[718]), .S(n4594), .Y(n3653) );
  MUX2X1 U4171 ( .B(fifo_array[616]), .A(fifo_array[650]), .S(n4594), .Y(n3657) );
  MUX2X1 U4172 ( .B(fifo_array[548]), .A(fifo_array[582]), .S(n4594), .Y(n3656) );
  MUX2X1 U4173 ( .B(n3655), .A(n3652), .S(n4655), .Y(n3659) );
  MUX2X1 U4174 ( .B(fifo_array[480]), .A(fifo_array[514]), .S(n4594), .Y(n3663) );
  MUX2X1 U4175 ( .B(fifo_array[412]), .A(fifo_array[446]), .S(n4594), .Y(n3662) );
  MUX2X1 U4176 ( .B(fifo_array[344]), .A(fifo_array[378]), .S(n4594), .Y(n3666) );
  MUX2X1 U4177 ( .B(fifo_array[276]), .A(fifo_array[310]), .S(n4594), .Y(n3665) );
  MUX2X1 U4178 ( .B(n3664), .A(n3661), .S(n4655), .Y(n3675) );
  MUX2X1 U4179 ( .B(fifo_array[208]), .A(fifo_array[242]), .S(n4595), .Y(n3669) );
  MUX2X1 U4180 ( .B(fifo_array[140]), .A(fifo_array[174]), .S(n4595), .Y(n3668) );
  MUX2X1 U4181 ( .B(fifo_array[72]), .A(fifo_array[106]), .S(n4595), .Y(n3672)
         );
  MUX2X1 U4182 ( .B(fifo_array[4]), .A(fifo_array[38]), .S(n4595), .Y(n3671)
         );
  MUX2X1 U4183 ( .B(n3670), .A(n3667), .S(n4655), .Y(n3674) );
  MUX2X1 U4184 ( .B(n3673), .A(n3658), .S(n23), .Y(n4550) );
  MUX2X1 U4185 ( .B(fifo_array[1025]), .A(fifo_array[1059]), .S(n4595), .Y(
        n3678) );
  MUX2X1 U4186 ( .B(fifo_array[957]), .A(fifo_array[991]), .S(n4595), .Y(n3677) );
  MUX2X1 U4187 ( .B(fifo_array[889]), .A(fifo_array[923]), .S(n4595), .Y(n3681) );
  MUX2X1 U4188 ( .B(fifo_array[821]), .A(fifo_array[855]), .S(n4595), .Y(n3680) );
  MUX2X1 U4189 ( .B(n3679), .A(n3676), .S(n4655), .Y(n3690) );
  MUX2X1 U4190 ( .B(fifo_array[753]), .A(fifo_array[787]), .S(n4595), .Y(n3684) );
  MUX2X1 U4191 ( .B(fifo_array[685]), .A(fifo_array[719]), .S(n4595), .Y(n3683) );
  MUX2X1 U4192 ( .B(fifo_array[617]), .A(fifo_array[651]), .S(n4595), .Y(n3687) );
  MUX2X1 U4193 ( .B(fifo_array[549]), .A(fifo_array[583]), .S(n4595), .Y(n3686) );
  MUX2X1 U4194 ( .B(n3685), .A(n3682), .S(n4655), .Y(n3689) );
  MUX2X1 U4195 ( .B(fifo_array[481]), .A(fifo_array[515]), .S(n4596), .Y(n3693) );
  MUX2X1 U4196 ( .B(fifo_array[413]), .A(fifo_array[447]), .S(n4596), .Y(n3692) );
  MUX2X1 U4197 ( .B(fifo_array[345]), .A(fifo_array[379]), .S(n4596), .Y(n3696) );
  MUX2X1 U4198 ( .B(fifo_array[277]), .A(fifo_array[311]), .S(n4596), .Y(n3695) );
  MUX2X1 U4199 ( .B(n3694), .A(n3691), .S(n4655), .Y(n3705) );
  MUX2X1 U4200 ( .B(fifo_array[209]), .A(fifo_array[243]), .S(n4596), .Y(n3699) );
  MUX2X1 U4201 ( .B(fifo_array[141]), .A(fifo_array[175]), .S(n4596), .Y(n3698) );
  MUX2X1 U4202 ( .B(fifo_array[73]), .A(fifo_array[107]), .S(n4596), .Y(n3702)
         );
  MUX2X1 U4203 ( .B(fifo_array[5]), .A(fifo_array[39]), .S(n4596), .Y(n3701)
         );
  MUX2X1 U4204 ( .B(n3700), .A(n3697), .S(n4655), .Y(n3704) );
  MUX2X1 U4205 ( .B(n3703), .A(n3688), .S(n23), .Y(n4551) );
  MUX2X1 U4206 ( .B(fifo_array[1026]), .A(fifo_array[1060]), .S(n4596), .Y(
        n3708) );
  MUX2X1 U4207 ( .B(fifo_array[958]), .A(fifo_array[992]), .S(n4596), .Y(n3707) );
  MUX2X1 U4208 ( .B(fifo_array[890]), .A(fifo_array[924]), .S(n4596), .Y(n3711) );
  MUX2X1 U4209 ( .B(fifo_array[822]), .A(fifo_array[856]), .S(n4596), .Y(n3710) );
  MUX2X1 U4210 ( .B(n3709), .A(n3706), .S(n4655), .Y(n3720) );
  MUX2X1 U4211 ( .B(fifo_array[754]), .A(fifo_array[788]), .S(n4597), .Y(n3714) );
  MUX2X1 U4212 ( .B(fifo_array[686]), .A(fifo_array[720]), .S(n4597), .Y(n3713) );
  MUX2X1 U4213 ( .B(fifo_array[618]), .A(fifo_array[652]), .S(n4597), .Y(n3717) );
  MUX2X1 U4214 ( .B(fifo_array[550]), .A(fifo_array[584]), .S(n4597), .Y(n3716) );
  MUX2X1 U4215 ( .B(n3715), .A(n3712), .S(n4655), .Y(n3719) );
  MUX2X1 U4216 ( .B(fifo_array[482]), .A(fifo_array[516]), .S(n4597), .Y(n3723) );
  MUX2X1 U4217 ( .B(fifo_array[414]), .A(fifo_array[448]), .S(n4597), .Y(n3722) );
  MUX2X1 U4218 ( .B(fifo_array[346]), .A(fifo_array[380]), .S(n4597), .Y(n3726) );
  MUX2X1 U4219 ( .B(fifo_array[278]), .A(fifo_array[312]), .S(n4597), .Y(n3725) );
  MUX2X1 U4220 ( .B(n3724), .A(n3721), .S(n4655), .Y(n3735) );
  MUX2X1 U4221 ( .B(fifo_array[210]), .A(fifo_array[244]), .S(n4597), .Y(n3729) );
  MUX2X1 U4222 ( .B(fifo_array[142]), .A(fifo_array[176]), .S(n4597), .Y(n3728) );
  MUX2X1 U4223 ( .B(fifo_array[74]), .A(fifo_array[108]), .S(n4597), .Y(n3732)
         );
  MUX2X1 U4224 ( .B(fifo_array[6]), .A(fifo_array[40]), .S(n4597), .Y(n3731)
         );
  MUX2X1 U4225 ( .B(n3730), .A(n3727), .S(n4655), .Y(n3734) );
  MUX2X1 U4226 ( .B(n3733), .A(n3718), .S(n23), .Y(n4552) );
  MUX2X1 U4227 ( .B(fifo_array[1027]), .A(fifo_array[1061]), .S(n4598), .Y(
        n3738) );
  MUX2X1 U4228 ( .B(fifo_array[959]), .A(fifo_array[993]), .S(n4598), .Y(n3737) );
  MUX2X1 U4229 ( .B(fifo_array[891]), .A(fifo_array[925]), .S(n4598), .Y(n3741) );
  MUX2X1 U4230 ( .B(fifo_array[823]), .A(fifo_array[857]), .S(n4598), .Y(n3740) );
  MUX2X1 U4231 ( .B(n3739), .A(n3736), .S(n21), .Y(n3750) );
  MUX2X1 U4232 ( .B(fifo_array[755]), .A(fifo_array[789]), .S(n4598), .Y(n3744) );
  MUX2X1 U4233 ( .B(fifo_array[687]), .A(fifo_array[721]), .S(n4598), .Y(n3743) );
  MUX2X1 U4234 ( .B(fifo_array[619]), .A(fifo_array[653]), .S(n4598), .Y(n3747) );
  MUX2X1 U4235 ( .B(fifo_array[551]), .A(fifo_array[585]), .S(n4598), .Y(n3746) );
  MUX2X1 U4236 ( .B(n3745), .A(n3742), .S(n21), .Y(n3749) );
  MUX2X1 U4237 ( .B(fifo_array[483]), .A(fifo_array[517]), .S(n4598), .Y(n3753) );
  MUX2X1 U4238 ( .B(fifo_array[415]), .A(fifo_array[449]), .S(n4598), .Y(n3752) );
  MUX2X1 U4239 ( .B(fifo_array[347]), .A(fifo_array[381]), .S(n4598), .Y(n3756) );
  MUX2X1 U4240 ( .B(fifo_array[279]), .A(fifo_array[313]), .S(n4598), .Y(n3755) );
  MUX2X1 U4241 ( .B(n3754), .A(n3751), .S(n21), .Y(n3765) );
  MUX2X1 U4242 ( .B(fifo_array[211]), .A(fifo_array[245]), .S(n4599), .Y(n3759) );
  MUX2X1 U4243 ( .B(fifo_array[143]), .A(fifo_array[177]), .S(n4599), .Y(n3758) );
  MUX2X1 U4244 ( .B(fifo_array[75]), .A(fifo_array[109]), .S(n4599), .Y(n3762)
         );
  MUX2X1 U4245 ( .B(fifo_array[7]), .A(fifo_array[41]), .S(n4599), .Y(n3761)
         );
  MUX2X1 U4246 ( .B(n3760), .A(n3757), .S(n21), .Y(n3764) );
  MUX2X1 U4247 ( .B(n3763), .A(n3748), .S(n23), .Y(n4553) );
  MUX2X1 U4248 ( .B(fifo_array[1028]), .A(fifo_array[1062]), .S(n4599), .Y(
        n3768) );
  MUX2X1 U4249 ( .B(fifo_array[960]), .A(fifo_array[994]), .S(n4599), .Y(n3767) );
  MUX2X1 U4250 ( .B(fifo_array[892]), .A(fifo_array[926]), .S(n4599), .Y(n3771) );
  MUX2X1 U4251 ( .B(fifo_array[824]), .A(fifo_array[858]), .S(n4599), .Y(n3770) );
  MUX2X1 U4252 ( .B(n3769), .A(n3766), .S(n21), .Y(n3780) );
  MUX2X1 U4253 ( .B(fifo_array[756]), .A(fifo_array[790]), .S(n4599), .Y(n3774) );
  MUX2X1 U4254 ( .B(fifo_array[688]), .A(fifo_array[722]), .S(n4599), .Y(n3773) );
  MUX2X1 U4255 ( .B(fifo_array[620]), .A(fifo_array[654]), .S(n4599), .Y(n3777) );
  MUX2X1 U4256 ( .B(fifo_array[552]), .A(fifo_array[586]), .S(n4599), .Y(n3776) );
  MUX2X1 U4257 ( .B(n3775), .A(n3772), .S(n21), .Y(n3779) );
  MUX2X1 U4258 ( .B(fifo_array[484]), .A(fifo_array[518]), .S(n4600), .Y(n3783) );
  MUX2X1 U4259 ( .B(fifo_array[416]), .A(fifo_array[450]), .S(n4600), .Y(n3782) );
  MUX2X1 U4260 ( .B(fifo_array[348]), .A(fifo_array[382]), .S(n4600), .Y(n3786) );
  MUX2X1 U4261 ( .B(fifo_array[280]), .A(fifo_array[314]), .S(n4600), .Y(n3785) );
  MUX2X1 U4262 ( .B(n3784), .A(n3781), .S(n21), .Y(n3795) );
  MUX2X1 U4263 ( .B(fifo_array[212]), .A(fifo_array[246]), .S(n4600), .Y(n3789) );
  MUX2X1 U4264 ( .B(fifo_array[144]), .A(fifo_array[178]), .S(n4600), .Y(n3788) );
  MUX2X1 U4265 ( .B(fifo_array[76]), .A(fifo_array[110]), .S(n4600), .Y(n3792)
         );
  MUX2X1 U4266 ( .B(fifo_array[8]), .A(fifo_array[42]), .S(n4600), .Y(n3791)
         );
  MUX2X1 U4267 ( .B(n3790), .A(n3787), .S(n21), .Y(n3794) );
  MUX2X1 U4268 ( .B(n3793), .A(n3778), .S(n23), .Y(n4554) );
  MUX2X1 U4269 ( .B(fifo_array[1029]), .A(fifo_array[1063]), .S(n4600), .Y(
        n3798) );
  MUX2X1 U4270 ( .B(fifo_array[961]), .A(fifo_array[995]), .S(n4600), .Y(n3797) );
  MUX2X1 U4271 ( .B(fifo_array[893]), .A(fifo_array[927]), .S(n4600), .Y(n3801) );
  MUX2X1 U4272 ( .B(fifo_array[825]), .A(fifo_array[859]), .S(n4600), .Y(n3800) );
  MUX2X1 U4273 ( .B(n3799), .A(n3796), .S(n21), .Y(n3810) );
  MUX2X1 U4274 ( .B(fifo_array[757]), .A(fifo_array[791]), .S(n4601), .Y(n3804) );
  MUX2X1 U4275 ( .B(fifo_array[689]), .A(fifo_array[723]), .S(n4601), .Y(n3803) );
  MUX2X1 U4276 ( .B(fifo_array[621]), .A(fifo_array[655]), .S(n4601), .Y(n3807) );
  MUX2X1 U4277 ( .B(fifo_array[553]), .A(fifo_array[587]), .S(n4601), .Y(n3806) );
  MUX2X1 U4278 ( .B(n3805), .A(n3802), .S(n21), .Y(n3809) );
  MUX2X1 U4279 ( .B(fifo_array[485]), .A(fifo_array[519]), .S(n4601), .Y(n3813) );
  MUX2X1 U4280 ( .B(fifo_array[417]), .A(fifo_array[451]), .S(n4601), .Y(n3812) );
  MUX2X1 U4281 ( .B(fifo_array[349]), .A(fifo_array[383]), .S(n4601), .Y(n3816) );
  MUX2X1 U4282 ( .B(fifo_array[281]), .A(fifo_array[315]), .S(n4601), .Y(n3815) );
  MUX2X1 U4283 ( .B(n3814), .A(n3811), .S(n21), .Y(n3825) );
  MUX2X1 U4284 ( .B(fifo_array[213]), .A(fifo_array[247]), .S(n4601), .Y(n3819) );
  MUX2X1 U4285 ( .B(fifo_array[145]), .A(fifo_array[179]), .S(n4601), .Y(n3818) );
  MUX2X1 U4286 ( .B(fifo_array[77]), .A(fifo_array[111]), .S(n4601), .Y(n3822)
         );
  MUX2X1 U4287 ( .B(fifo_array[9]), .A(fifo_array[43]), .S(n4601), .Y(n3821)
         );
  MUX2X1 U4288 ( .B(n3820), .A(n3817), .S(n21), .Y(n3824) );
  MUX2X1 U4289 ( .B(n3823), .A(n3808), .S(n23), .Y(n4555) );
  MUX2X1 U4290 ( .B(fifo_array[1030]), .A(fifo_array[1064]), .S(n4602), .Y(
        n3828) );
  MUX2X1 U4291 ( .B(fifo_array[962]), .A(fifo_array[996]), .S(n4602), .Y(n3827) );
  MUX2X1 U4292 ( .B(fifo_array[894]), .A(fifo_array[928]), .S(n4602), .Y(n3831) );
  MUX2X1 U4293 ( .B(fifo_array[826]), .A(fifo_array[860]), .S(n4602), .Y(n3830) );
  MUX2X1 U4294 ( .B(n3829), .A(n3826), .S(n21), .Y(n3840) );
  MUX2X1 U4295 ( .B(fifo_array[758]), .A(fifo_array[792]), .S(n4602), .Y(n3834) );
  MUX2X1 U4296 ( .B(fifo_array[690]), .A(fifo_array[724]), .S(n4602), .Y(n3833) );
  MUX2X1 U4297 ( .B(fifo_array[622]), .A(fifo_array[656]), .S(n4602), .Y(n3837) );
  MUX2X1 U4298 ( .B(fifo_array[554]), .A(fifo_array[588]), .S(n4602), .Y(n3836) );
  MUX2X1 U4299 ( .B(n3835), .A(n3832), .S(n21), .Y(n3839) );
  MUX2X1 U4300 ( .B(fifo_array[486]), .A(fifo_array[520]), .S(n4602), .Y(n3843) );
  MUX2X1 U4301 ( .B(fifo_array[418]), .A(fifo_array[452]), .S(n4602), .Y(n3842) );
  MUX2X1 U4302 ( .B(fifo_array[350]), .A(fifo_array[384]), .S(n4602), .Y(n3846) );
  MUX2X1 U4303 ( .B(fifo_array[282]), .A(fifo_array[316]), .S(n4602), .Y(n3845) );
  MUX2X1 U4304 ( .B(n3844), .A(n3841), .S(n21), .Y(n3855) );
  MUX2X1 U4305 ( .B(fifo_array[214]), .A(fifo_array[248]), .S(n4603), .Y(n3849) );
  MUX2X1 U4306 ( .B(fifo_array[146]), .A(fifo_array[180]), .S(n4603), .Y(n3848) );
  MUX2X1 U4307 ( .B(fifo_array[78]), .A(fifo_array[112]), .S(n4603), .Y(n3852)
         );
  MUX2X1 U4308 ( .B(fifo_array[10]), .A(fifo_array[44]), .S(n4603), .Y(n3851)
         );
  MUX2X1 U4309 ( .B(n3850), .A(n3847), .S(n21), .Y(n3854) );
  MUX2X1 U4310 ( .B(n3853), .A(n3838), .S(n23), .Y(n4556) );
  MUX2X1 U4311 ( .B(fifo_array[1031]), .A(fifo_array[1065]), .S(n4603), .Y(
        n3858) );
  MUX2X1 U4312 ( .B(fifo_array[963]), .A(fifo_array[997]), .S(n4603), .Y(n3857) );
  MUX2X1 U4313 ( .B(fifo_array[895]), .A(fifo_array[929]), .S(n4603), .Y(n3861) );
  MUX2X1 U4314 ( .B(fifo_array[827]), .A(fifo_array[861]), .S(n4603), .Y(n3860) );
  MUX2X1 U4315 ( .B(n3859), .A(n3856), .S(n21), .Y(n3870) );
  MUX2X1 U4316 ( .B(fifo_array[759]), .A(fifo_array[793]), .S(n4603), .Y(n3864) );
  MUX2X1 U4317 ( .B(fifo_array[691]), .A(fifo_array[725]), .S(n4603), .Y(n3863) );
  MUX2X1 U4318 ( .B(fifo_array[623]), .A(fifo_array[657]), .S(n4603), .Y(n3867) );
  MUX2X1 U4319 ( .B(fifo_array[555]), .A(fifo_array[589]), .S(n4603), .Y(n3866) );
  MUX2X1 U4320 ( .B(n3865), .A(n3862), .S(n21), .Y(n3869) );
  MUX2X1 U4321 ( .B(fifo_array[487]), .A(fifo_array[521]), .S(n4604), .Y(n3873) );
  MUX2X1 U4322 ( .B(fifo_array[419]), .A(fifo_array[453]), .S(n4604), .Y(n3872) );
  MUX2X1 U4323 ( .B(fifo_array[351]), .A(fifo_array[385]), .S(n4604), .Y(n3876) );
  MUX2X1 U4324 ( .B(fifo_array[283]), .A(fifo_array[317]), .S(n4604), .Y(n3875) );
  MUX2X1 U4325 ( .B(n3874), .A(n3871), .S(n21), .Y(n3885) );
  MUX2X1 U4326 ( .B(fifo_array[215]), .A(fifo_array[249]), .S(n4604), .Y(n3879) );
  MUX2X1 U4327 ( .B(fifo_array[147]), .A(fifo_array[181]), .S(n4604), .Y(n3878) );
  MUX2X1 U4328 ( .B(fifo_array[79]), .A(fifo_array[113]), .S(n4604), .Y(n3882)
         );
  MUX2X1 U4329 ( .B(fifo_array[11]), .A(fifo_array[45]), .S(n4604), .Y(n3881)
         );
  MUX2X1 U4330 ( .B(n3880), .A(n3877), .S(n21), .Y(n3884) );
  MUX2X1 U4331 ( .B(n3883), .A(n3868), .S(n23), .Y(n4557) );
  MUX2X1 U4332 ( .B(fifo_array[1032]), .A(fifo_array[1066]), .S(n4604), .Y(
        n3888) );
  MUX2X1 U4333 ( .B(fifo_array[964]), .A(fifo_array[998]), .S(n4604), .Y(n3887) );
  MUX2X1 U4334 ( .B(fifo_array[896]), .A(fifo_array[930]), .S(n4604), .Y(n3891) );
  MUX2X1 U4335 ( .B(fifo_array[828]), .A(fifo_array[862]), .S(n4604), .Y(n3890) );
  MUX2X1 U4336 ( .B(n3889), .A(n3886), .S(n21), .Y(n3900) );
  MUX2X1 U4337 ( .B(fifo_array[760]), .A(fifo_array[794]), .S(n4605), .Y(n3894) );
  MUX2X1 U4338 ( .B(fifo_array[692]), .A(fifo_array[726]), .S(n4605), .Y(n3893) );
  MUX2X1 U4339 ( .B(fifo_array[624]), .A(fifo_array[658]), .S(n4605), .Y(n3897) );
  MUX2X1 U4340 ( .B(fifo_array[556]), .A(fifo_array[590]), .S(n4605), .Y(n3896) );
  MUX2X1 U4341 ( .B(n3895), .A(n3892), .S(n21), .Y(n3899) );
  MUX2X1 U4342 ( .B(fifo_array[488]), .A(fifo_array[522]), .S(n4605), .Y(n3903) );
  MUX2X1 U4343 ( .B(fifo_array[420]), .A(fifo_array[454]), .S(n4605), .Y(n3902) );
  MUX2X1 U4344 ( .B(fifo_array[352]), .A(fifo_array[386]), .S(n4605), .Y(n3906) );
  MUX2X1 U4345 ( .B(fifo_array[284]), .A(fifo_array[318]), .S(n4605), .Y(n3905) );
  MUX2X1 U4346 ( .B(n3904), .A(n3901), .S(n21), .Y(n3915) );
  MUX2X1 U4347 ( .B(fifo_array[216]), .A(fifo_array[250]), .S(n4605), .Y(n3909) );
  MUX2X1 U4348 ( .B(fifo_array[148]), .A(fifo_array[182]), .S(n4605), .Y(n3908) );
  MUX2X1 U4349 ( .B(fifo_array[80]), .A(fifo_array[114]), .S(n4605), .Y(n3912)
         );
  MUX2X1 U4350 ( .B(fifo_array[12]), .A(fifo_array[46]), .S(n4605), .Y(n3911)
         );
  MUX2X1 U4351 ( .B(n3910), .A(n3907), .S(n21), .Y(n3914) );
  MUX2X1 U4352 ( .B(n3913), .A(n3898), .S(n23), .Y(n4558) );
  MUX2X1 U4353 ( .B(fifo_array[1033]), .A(fifo_array[1067]), .S(n4606), .Y(
        n3918) );
  MUX2X1 U4354 ( .B(fifo_array[965]), .A(fifo_array[999]), .S(n4606), .Y(n3917) );
  MUX2X1 U4355 ( .B(fifo_array[897]), .A(fifo_array[931]), .S(n4606), .Y(n3921) );
  MUX2X1 U4356 ( .B(fifo_array[829]), .A(fifo_array[863]), .S(n4606), .Y(n3920) );
  MUX2X1 U4357 ( .B(n3919), .A(n3916), .S(n21), .Y(n3930) );
  MUX2X1 U4358 ( .B(fifo_array[761]), .A(fifo_array[795]), .S(n4606), .Y(n3924) );
  MUX2X1 U4359 ( .B(fifo_array[693]), .A(fifo_array[727]), .S(n4606), .Y(n3923) );
  MUX2X1 U4360 ( .B(fifo_array[625]), .A(fifo_array[659]), .S(n4606), .Y(n3927) );
  MUX2X1 U4361 ( .B(fifo_array[557]), .A(fifo_array[591]), .S(n4606), .Y(n3926) );
  MUX2X1 U4362 ( .B(n3925), .A(n3922), .S(n21), .Y(n3929) );
  MUX2X1 U4363 ( .B(fifo_array[489]), .A(fifo_array[523]), .S(n4606), .Y(n3933) );
  MUX2X1 U4364 ( .B(fifo_array[421]), .A(fifo_array[455]), .S(n4606), .Y(n3932) );
  MUX2X1 U4365 ( .B(fifo_array[353]), .A(fifo_array[387]), .S(n4606), .Y(n3936) );
  MUX2X1 U4366 ( .B(fifo_array[285]), .A(fifo_array[319]), .S(n4606), .Y(n3935) );
  MUX2X1 U4367 ( .B(n3934), .A(n3931), .S(n21), .Y(n3945) );
  MUX2X1 U4368 ( .B(fifo_array[217]), .A(fifo_array[251]), .S(n4607), .Y(n3939) );
  MUX2X1 U4369 ( .B(fifo_array[149]), .A(fifo_array[183]), .S(n4607), .Y(n3938) );
  MUX2X1 U4370 ( .B(fifo_array[81]), .A(fifo_array[115]), .S(n4607), .Y(n3942)
         );
  MUX2X1 U4371 ( .B(fifo_array[13]), .A(fifo_array[47]), .S(n4607), .Y(n3941)
         );
  MUX2X1 U4372 ( .B(n3940), .A(n3937), .S(n21), .Y(n3944) );
  MUX2X1 U4373 ( .B(n3943), .A(n3928), .S(n23), .Y(n4559) );
  MUX2X1 U4374 ( .B(fifo_array[1034]), .A(fifo_array[1068]), .S(n4607), .Y(
        n3948) );
  MUX2X1 U4375 ( .B(fifo_array[966]), .A(fifo_array[1000]), .S(n4607), .Y(
        n3947) );
  MUX2X1 U4376 ( .B(fifo_array[898]), .A(fifo_array[932]), .S(n4607), .Y(n3951) );
  MUX2X1 U4377 ( .B(fifo_array[830]), .A(fifo_array[864]), .S(n4607), .Y(n3950) );
  MUX2X1 U4378 ( .B(n3949), .A(n3946), .S(n21), .Y(n3960) );
  MUX2X1 U4379 ( .B(fifo_array[762]), .A(fifo_array[796]), .S(n4607), .Y(n3954) );
  MUX2X1 U4380 ( .B(fifo_array[694]), .A(fifo_array[728]), .S(n4607), .Y(n3953) );
  MUX2X1 U4381 ( .B(fifo_array[626]), .A(fifo_array[660]), .S(n4607), .Y(n3957) );
  MUX2X1 U4382 ( .B(fifo_array[558]), .A(fifo_array[592]), .S(n4607), .Y(n3956) );
  MUX2X1 U4383 ( .B(n3955), .A(n3952), .S(n21), .Y(n3959) );
  MUX2X1 U4384 ( .B(fifo_array[490]), .A(fifo_array[524]), .S(n4608), .Y(n3963) );
  MUX2X1 U4385 ( .B(fifo_array[422]), .A(fifo_array[456]), .S(n4608), .Y(n3962) );
  MUX2X1 U4386 ( .B(fifo_array[354]), .A(fifo_array[388]), .S(n4608), .Y(n3966) );
  MUX2X1 U4387 ( .B(fifo_array[286]), .A(fifo_array[320]), .S(n4608), .Y(n3965) );
  MUX2X1 U4388 ( .B(n3964), .A(n3961), .S(n21), .Y(n3975) );
  MUX2X1 U4389 ( .B(fifo_array[218]), .A(fifo_array[252]), .S(n4608), .Y(n3969) );
  MUX2X1 U4390 ( .B(fifo_array[150]), .A(fifo_array[184]), .S(n4608), .Y(n3968) );
  MUX2X1 U4391 ( .B(fifo_array[82]), .A(fifo_array[116]), .S(n4608), .Y(n3972)
         );
  MUX2X1 U4392 ( .B(fifo_array[14]), .A(fifo_array[48]), .S(n4608), .Y(n3971)
         );
  MUX2X1 U4393 ( .B(n3970), .A(n3967), .S(n21), .Y(n3974) );
  MUX2X1 U4394 ( .B(n3973), .A(n3958), .S(n23), .Y(n4560) );
  MUX2X1 U4395 ( .B(fifo_array[1035]), .A(fifo_array[1069]), .S(n4608), .Y(
        n3978) );
  MUX2X1 U4396 ( .B(fifo_array[967]), .A(fifo_array[1001]), .S(n4608), .Y(
        n3977) );
  MUX2X1 U4397 ( .B(fifo_array[899]), .A(fifo_array[933]), .S(n4608), .Y(n3981) );
  MUX2X1 U4398 ( .B(fifo_array[831]), .A(fifo_array[865]), .S(n4608), .Y(n3980) );
  MUX2X1 U4399 ( .B(n3979), .A(n3976), .S(n21), .Y(n3990) );
  MUX2X1 U4400 ( .B(fifo_array[763]), .A(fifo_array[797]), .S(n4609), .Y(n3984) );
  MUX2X1 U4401 ( .B(fifo_array[695]), .A(fifo_array[729]), .S(n4609), .Y(n3983) );
  MUX2X1 U4402 ( .B(fifo_array[627]), .A(fifo_array[661]), .S(n4609), .Y(n3987) );
  MUX2X1 U4403 ( .B(fifo_array[559]), .A(fifo_array[593]), .S(n4609), .Y(n3986) );
  MUX2X1 U4404 ( .B(n3985), .A(n3982), .S(n21), .Y(n3989) );
  MUX2X1 U4405 ( .B(fifo_array[491]), .A(fifo_array[525]), .S(n4609), .Y(n3993) );
  MUX2X1 U4406 ( .B(fifo_array[423]), .A(fifo_array[457]), .S(n4609), .Y(n3992) );
  MUX2X1 U4407 ( .B(fifo_array[355]), .A(fifo_array[389]), .S(n4609), .Y(n3996) );
  MUX2X1 U4408 ( .B(fifo_array[287]), .A(fifo_array[321]), .S(n4609), .Y(n3995) );
  MUX2X1 U4409 ( .B(n3994), .A(n3991), .S(n21), .Y(n4005) );
  MUX2X1 U4410 ( .B(fifo_array[219]), .A(fifo_array[253]), .S(n4609), .Y(n3999) );
  MUX2X1 U4411 ( .B(fifo_array[151]), .A(fifo_array[185]), .S(n4609), .Y(n3998) );
  MUX2X1 U4412 ( .B(fifo_array[83]), .A(fifo_array[117]), .S(n4609), .Y(n4002)
         );
  MUX2X1 U4413 ( .B(fifo_array[15]), .A(fifo_array[49]), .S(n4609), .Y(n4001)
         );
  MUX2X1 U4414 ( .B(n4000), .A(n3997), .S(n21), .Y(n4004) );
  MUX2X1 U4415 ( .B(n4003), .A(n3988), .S(n23), .Y(n4561) );
  MUX2X1 U4416 ( .B(fifo_array[1036]), .A(fifo_array[1070]), .S(n4610), .Y(
        n4008) );
  MUX2X1 U4417 ( .B(fifo_array[968]), .A(fifo_array[1002]), .S(n4610), .Y(
        n4007) );
  MUX2X1 U4418 ( .B(fifo_array[900]), .A(fifo_array[934]), .S(n4610), .Y(n4011) );
  MUX2X1 U4419 ( .B(fifo_array[832]), .A(fifo_array[866]), .S(n4610), .Y(n4010) );
  MUX2X1 U4420 ( .B(n4009), .A(n4006), .S(n21), .Y(n4020) );
  MUX2X1 U4421 ( .B(fifo_array[764]), .A(fifo_array[798]), .S(n4610), .Y(n4014) );
  MUX2X1 U4422 ( .B(fifo_array[696]), .A(fifo_array[730]), .S(n4610), .Y(n4013) );
  MUX2X1 U4423 ( .B(fifo_array[628]), .A(fifo_array[662]), .S(n4610), .Y(n4017) );
  MUX2X1 U4424 ( .B(fifo_array[560]), .A(fifo_array[594]), .S(n4610), .Y(n4016) );
  MUX2X1 U4425 ( .B(n4015), .A(n4012), .S(n21), .Y(n4019) );
  MUX2X1 U4426 ( .B(fifo_array[492]), .A(fifo_array[526]), .S(n4610), .Y(n4023) );
  MUX2X1 U4427 ( .B(fifo_array[424]), .A(fifo_array[458]), .S(n4610), .Y(n4022) );
  MUX2X1 U4428 ( .B(fifo_array[356]), .A(fifo_array[390]), .S(n4610), .Y(n4026) );
  MUX2X1 U4429 ( .B(fifo_array[288]), .A(fifo_array[322]), .S(n4610), .Y(n4025) );
  MUX2X1 U4430 ( .B(n4024), .A(n4021), .S(n21), .Y(n4035) );
  MUX2X1 U4431 ( .B(fifo_array[220]), .A(fifo_array[254]), .S(n4611), .Y(n4029) );
  MUX2X1 U4432 ( .B(fifo_array[152]), .A(fifo_array[186]), .S(n4611), .Y(n4028) );
  MUX2X1 U4433 ( .B(fifo_array[84]), .A(fifo_array[118]), .S(n4611), .Y(n4032)
         );
  MUX2X1 U4434 ( .B(fifo_array[16]), .A(fifo_array[50]), .S(n4611), .Y(n4031)
         );
  MUX2X1 U4435 ( .B(n4030), .A(n4027), .S(n21), .Y(n4034) );
  MUX2X1 U4436 ( .B(n4033), .A(n4018), .S(n23), .Y(n4562) );
  MUX2X1 U4437 ( .B(fifo_array[1037]), .A(fifo_array[1071]), .S(n4611), .Y(
        n4038) );
  MUX2X1 U4438 ( .B(fifo_array[969]), .A(fifo_array[1003]), .S(n4611), .Y(
        n4037) );
  MUX2X1 U4439 ( .B(fifo_array[901]), .A(fifo_array[935]), .S(n4611), .Y(n4041) );
  MUX2X1 U4440 ( .B(fifo_array[833]), .A(fifo_array[867]), .S(n4611), .Y(n4040) );
  MUX2X1 U4441 ( .B(n4039), .A(n4036), .S(n21), .Y(n4050) );
  MUX2X1 U4442 ( .B(fifo_array[765]), .A(fifo_array[799]), .S(n4611), .Y(n4044) );
  MUX2X1 U4443 ( .B(fifo_array[697]), .A(fifo_array[731]), .S(n4611), .Y(n4043) );
  MUX2X1 U4444 ( .B(fifo_array[629]), .A(fifo_array[663]), .S(n4611), .Y(n4047) );
  MUX2X1 U4445 ( .B(fifo_array[561]), .A(fifo_array[595]), .S(n4611), .Y(n4046) );
  MUX2X1 U4446 ( .B(n4045), .A(n4042), .S(n21), .Y(n4049) );
  MUX2X1 U4447 ( .B(fifo_array[493]), .A(fifo_array[527]), .S(n4612), .Y(n4053) );
  MUX2X1 U4448 ( .B(fifo_array[425]), .A(fifo_array[459]), .S(n4612), .Y(n4052) );
  MUX2X1 U4449 ( .B(fifo_array[357]), .A(fifo_array[391]), .S(n4612), .Y(n4056) );
  MUX2X1 U4450 ( .B(fifo_array[289]), .A(fifo_array[323]), .S(n4612), .Y(n4055) );
  MUX2X1 U4451 ( .B(n4054), .A(n4051), .S(n21), .Y(n4065) );
  MUX2X1 U4452 ( .B(fifo_array[221]), .A(fifo_array[255]), .S(n4612), .Y(n4059) );
  MUX2X1 U4453 ( .B(fifo_array[153]), .A(fifo_array[187]), .S(n4612), .Y(n4058) );
  MUX2X1 U4454 ( .B(fifo_array[85]), .A(fifo_array[119]), .S(n4612), .Y(n4062)
         );
  MUX2X1 U4455 ( .B(fifo_array[17]), .A(fifo_array[51]), .S(n4612), .Y(n4061)
         );
  MUX2X1 U4456 ( .B(n4060), .A(n4057), .S(n21), .Y(n4064) );
  MUX2X1 U4457 ( .B(n4063), .A(n4048), .S(n23), .Y(n4563) );
  MUX2X1 U4458 ( .B(fifo_array[1038]), .A(fifo_array[1072]), .S(n4612), .Y(
        n4068) );
  MUX2X1 U4459 ( .B(fifo_array[970]), .A(fifo_array[1004]), .S(n4612), .Y(
        n4067) );
  MUX2X1 U4460 ( .B(fifo_array[902]), .A(fifo_array[936]), .S(n4612), .Y(n4071) );
  MUX2X1 U4461 ( .B(fifo_array[834]), .A(fifo_array[868]), .S(n4612), .Y(n4070) );
  MUX2X1 U4462 ( .B(n4069), .A(n4066), .S(n21), .Y(n4080) );
  MUX2X1 U4463 ( .B(fifo_array[766]), .A(fifo_array[800]), .S(n4613), .Y(n4074) );
  MUX2X1 U4464 ( .B(fifo_array[698]), .A(fifo_array[732]), .S(n4613), .Y(n4073) );
  MUX2X1 U4465 ( .B(fifo_array[630]), .A(fifo_array[664]), .S(n4613), .Y(n4077) );
  MUX2X1 U4466 ( .B(fifo_array[562]), .A(fifo_array[596]), .S(n4613), .Y(n4076) );
  MUX2X1 U4467 ( .B(n4075), .A(n4072), .S(n21), .Y(n4079) );
  MUX2X1 U4468 ( .B(fifo_array[494]), .A(fifo_array[528]), .S(n4613), .Y(n4083) );
  MUX2X1 U4469 ( .B(fifo_array[426]), .A(fifo_array[460]), .S(n4613), .Y(n4082) );
  MUX2X1 U4470 ( .B(fifo_array[358]), .A(fifo_array[392]), .S(n4613), .Y(n4086) );
  MUX2X1 U4471 ( .B(fifo_array[290]), .A(fifo_array[324]), .S(n4613), .Y(n4085) );
  MUX2X1 U4472 ( .B(n4084), .A(n4081), .S(n21), .Y(n4095) );
  MUX2X1 U4473 ( .B(fifo_array[222]), .A(fifo_array[256]), .S(n4613), .Y(n4089) );
  MUX2X1 U4474 ( .B(fifo_array[154]), .A(fifo_array[188]), .S(n4613), .Y(n4088) );
  MUX2X1 U4475 ( .B(fifo_array[86]), .A(fifo_array[120]), .S(n4613), .Y(n4092)
         );
  MUX2X1 U4476 ( .B(fifo_array[18]), .A(fifo_array[52]), .S(n4613), .Y(n4091)
         );
  MUX2X1 U4477 ( .B(n4090), .A(n4087), .S(n21), .Y(n4094) );
  MUX2X1 U4478 ( .B(n4093), .A(n4078), .S(n23), .Y(n4564) );
  MUX2X1 U4479 ( .B(fifo_array[1039]), .A(fifo_array[1073]), .S(n4614), .Y(
        n4098) );
  MUX2X1 U4480 ( .B(fifo_array[971]), .A(fifo_array[1005]), .S(n4614), .Y(
        n4097) );
  MUX2X1 U4481 ( .B(fifo_array[903]), .A(fifo_array[937]), .S(n4614), .Y(n4101) );
  MUX2X1 U4482 ( .B(fifo_array[835]), .A(fifo_array[869]), .S(n4614), .Y(n4100) );
  MUX2X1 U4483 ( .B(n4099), .A(n4096), .S(n21), .Y(n4110) );
  MUX2X1 U4484 ( .B(fifo_array[767]), .A(fifo_array[801]), .S(n4614), .Y(n4104) );
  MUX2X1 U4485 ( .B(fifo_array[699]), .A(fifo_array[733]), .S(n4614), .Y(n4103) );
  MUX2X1 U4486 ( .B(fifo_array[631]), .A(fifo_array[665]), .S(n4614), .Y(n4107) );
  MUX2X1 U4487 ( .B(fifo_array[563]), .A(fifo_array[597]), .S(n4614), .Y(n4106) );
  MUX2X1 U4488 ( .B(n4105), .A(n4102), .S(n21), .Y(n4109) );
  MUX2X1 U4489 ( .B(fifo_array[495]), .A(fifo_array[529]), .S(n4614), .Y(n4113) );
  MUX2X1 U4490 ( .B(fifo_array[427]), .A(fifo_array[461]), .S(n4614), .Y(n4112) );
  MUX2X1 U4491 ( .B(fifo_array[359]), .A(fifo_array[393]), .S(n4614), .Y(n4116) );
  MUX2X1 U4492 ( .B(fifo_array[291]), .A(fifo_array[325]), .S(n4614), .Y(n4115) );
  MUX2X1 U4493 ( .B(n4114), .A(n4111), .S(n21), .Y(n4125) );
  MUX2X1 U4494 ( .B(fifo_array[223]), .A(fifo_array[257]), .S(n4615), .Y(n4119) );
  MUX2X1 U4495 ( .B(fifo_array[155]), .A(fifo_array[189]), .S(n4615), .Y(n4118) );
  MUX2X1 U4496 ( .B(fifo_array[87]), .A(fifo_array[121]), .S(n4615), .Y(n4122)
         );
  MUX2X1 U4497 ( .B(fifo_array[19]), .A(fifo_array[53]), .S(n4615), .Y(n4121)
         );
  MUX2X1 U4498 ( .B(n4120), .A(n4117), .S(n21), .Y(n4124) );
  MUX2X1 U4499 ( .B(n4123), .A(n4108), .S(n23), .Y(n4565) );
  MUX2X1 U4500 ( .B(fifo_array[1040]), .A(fifo_array[1074]), .S(n4615), .Y(
        n4128) );
  MUX2X1 U4501 ( .B(fifo_array[972]), .A(fifo_array[1006]), .S(n4615), .Y(
        n4127) );
  MUX2X1 U4502 ( .B(fifo_array[904]), .A(fifo_array[938]), .S(n4615), .Y(n4131) );
  MUX2X1 U4503 ( .B(fifo_array[836]), .A(fifo_array[870]), .S(n4615), .Y(n4130) );
  MUX2X1 U4504 ( .B(n4129), .A(n4126), .S(n21), .Y(n4140) );
  MUX2X1 U4505 ( .B(fifo_array[768]), .A(fifo_array[802]), .S(n4615), .Y(n4134) );
  MUX2X1 U4506 ( .B(fifo_array[700]), .A(fifo_array[734]), .S(n4615), .Y(n4133) );
  MUX2X1 U4507 ( .B(fifo_array[632]), .A(fifo_array[666]), .S(n4615), .Y(n4137) );
  MUX2X1 U4508 ( .B(fifo_array[564]), .A(fifo_array[598]), .S(n4615), .Y(n4136) );
  MUX2X1 U4509 ( .B(n4135), .A(n4132), .S(n21), .Y(n4139) );
  MUX2X1 U4510 ( .B(fifo_array[496]), .A(fifo_array[530]), .S(n4616), .Y(n4143) );
  MUX2X1 U4511 ( .B(fifo_array[428]), .A(fifo_array[462]), .S(n4616), .Y(n4142) );
  MUX2X1 U4512 ( .B(fifo_array[360]), .A(fifo_array[394]), .S(n4616), .Y(n4146) );
  MUX2X1 U4513 ( .B(fifo_array[292]), .A(fifo_array[326]), .S(n4616), .Y(n4145) );
  MUX2X1 U4514 ( .B(n4144), .A(n4141), .S(n21), .Y(n4155) );
  MUX2X1 U4515 ( .B(fifo_array[224]), .A(fifo_array[258]), .S(n4616), .Y(n4149) );
  MUX2X1 U4516 ( .B(fifo_array[156]), .A(fifo_array[190]), .S(n4616), .Y(n4148) );
  MUX2X1 U4517 ( .B(fifo_array[88]), .A(fifo_array[122]), .S(n4616), .Y(n4152)
         );
  MUX2X1 U4518 ( .B(fifo_array[20]), .A(fifo_array[54]), .S(n4616), .Y(n4151)
         );
  MUX2X1 U4519 ( .B(n4150), .A(n4147), .S(n21), .Y(n4154) );
  MUX2X1 U4520 ( .B(n4153), .A(n4138), .S(n23), .Y(n4566) );
  MUX2X1 U4521 ( .B(fifo_array[1041]), .A(fifo_array[1075]), .S(n4616), .Y(
        n4158) );
  MUX2X1 U4522 ( .B(fifo_array[973]), .A(fifo_array[1007]), .S(n4616), .Y(
        n4157) );
  MUX2X1 U4523 ( .B(fifo_array[905]), .A(fifo_array[939]), .S(n4616), .Y(n4161) );
  MUX2X1 U4524 ( .B(fifo_array[837]), .A(fifo_array[871]), .S(n4616), .Y(n4160) );
  MUX2X1 U4525 ( .B(n4159), .A(n4156), .S(n21), .Y(n4170) );
  MUX2X1 U4526 ( .B(fifo_array[769]), .A(fifo_array[803]), .S(n4617), .Y(n4164) );
  MUX2X1 U4527 ( .B(fifo_array[701]), .A(fifo_array[735]), .S(n4617), .Y(n4163) );
  MUX2X1 U4528 ( .B(fifo_array[633]), .A(fifo_array[667]), .S(n4617), .Y(n4167) );
  MUX2X1 U4529 ( .B(fifo_array[565]), .A(fifo_array[599]), .S(n4617), .Y(n4166) );
  MUX2X1 U4530 ( .B(n4165), .A(n4162), .S(n21), .Y(n4169) );
  MUX2X1 U4531 ( .B(fifo_array[497]), .A(fifo_array[531]), .S(n4617), .Y(n4173) );
  MUX2X1 U4532 ( .B(fifo_array[429]), .A(fifo_array[463]), .S(n4617), .Y(n4172) );
  MUX2X1 U4533 ( .B(fifo_array[361]), .A(fifo_array[395]), .S(n4617), .Y(n4176) );
  MUX2X1 U4534 ( .B(fifo_array[293]), .A(fifo_array[327]), .S(n4617), .Y(n4175) );
  MUX2X1 U4535 ( .B(n4174), .A(n4171), .S(n21), .Y(n4185) );
  MUX2X1 U4536 ( .B(fifo_array[225]), .A(fifo_array[259]), .S(n4617), .Y(n4179) );
  MUX2X1 U4537 ( .B(fifo_array[157]), .A(fifo_array[191]), .S(n4617), .Y(n4178) );
  MUX2X1 U4538 ( .B(fifo_array[89]), .A(fifo_array[123]), .S(n4617), .Y(n4182)
         );
  MUX2X1 U4539 ( .B(fifo_array[21]), .A(fifo_array[55]), .S(n4617), .Y(n4181)
         );
  MUX2X1 U4540 ( .B(n4180), .A(n4177), .S(n21), .Y(n4184) );
  MUX2X1 U4541 ( .B(n4183), .A(n4168), .S(n23), .Y(n4567) );
  MUX2X1 U4542 ( .B(fifo_array[1042]), .A(fifo_array[1076]), .S(n4618), .Y(
        n4188) );
  MUX2X1 U4543 ( .B(fifo_array[974]), .A(fifo_array[1008]), .S(n4618), .Y(
        n4187) );
  MUX2X1 U4544 ( .B(fifo_array[906]), .A(fifo_array[940]), .S(n4618), .Y(n4191) );
  MUX2X1 U4545 ( .B(fifo_array[838]), .A(fifo_array[872]), .S(n4618), .Y(n4190) );
  MUX2X1 U4546 ( .B(n4189), .A(n4186), .S(n21), .Y(n4200) );
  MUX2X1 U4547 ( .B(fifo_array[770]), .A(fifo_array[804]), .S(n4618), .Y(n4194) );
  MUX2X1 U4548 ( .B(fifo_array[702]), .A(fifo_array[736]), .S(n4618), .Y(n4193) );
  MUX2X1 U4549 ( .B(fifo_array[634]), .A(fifo_array[668]), .S(n4618), .Y(n4197) );
  MUX2X1 U4550 ( .B(fifo_array[566]), .A(fifo_array[600]), .S(n4618), .Y(n4196) );
  MUX2X1 U4551 ( .B(n4195), .A(n4192), .S(n21), .Y(n4199) );
  MUX2X1 U4552 ( .B(fifo_array[498]), .A(fifo_array[532]), .S(n4618), .Y(n4203) );
  MUX2X1 U4553 ( .B(fifo_array[430]), .A(fifo_array[464]), .S(n4618), .Y(n4202) );
  MUX2X1 U4554 ( .B(fifo_array[362]), .A(fifo_array[396]), .S(n4618), .Y(n4206) );
  MUX2X1 U4555 ( .B(fifo_array[294]), .A(fifo_array[328]), .S(n4618), .Y(n4205) );
  MUX2X1 U4556 ( .B(n4204), .A(n4201), .S(n21), .Y(n4215) );
  MUX2X1 U4557 ( .B(fifo_array[226]), .A(fifo_array[260]), .S(n4619), .Y(n4209) );
  MUX2X1 U4558 ( .B(fifo_array[158]), .A(fifo_array[192]), .S(n4619), .Y(n4208) );
  MUX2X1 U4559 ( .B(fifo_array[90]), .A(fifo_array[124]), .S(n4619), .Y(n4212)
         );
  MUX2X1 U4560 ( .B(fifo_array[22]), .A(fifo_array[56]), .S(n4619), .Y(n4211)
         );
  MUX2X1 U4561 ( .B(n4210), .A(n4207), .S(n21), .Y(n4214) );
  MUX2X1 U4562 ( .B(n4213), .A(n4198), .S(n23), .Y(n4568) );
  MUX2X1 U4563 ( .B(fifo_array[1043]), .A(fifo_array[1077]), .S(n4619), .Y(
        n4218) );
  MUX2X1 U4564 ( .B(fifo_array[975]), .A(fifo_array[1009]), .S(n4619), .Y(
        n4217) );
  MUX2X1 U4565 ( .B(fifo_array[907]), .A(fifo_array[941]), .S(n4619), .Y(n4221) );
  MUX2X1 U4566 ( .B(fifo_array[839]), .A(fifo_array[873]), .S(n4619), .Y(n4220) );
  MUX2X1 U4567 ( .B(n4219), .A(n4216), .S(n4654), .Y(n4230) );
  MUX2X1 U4568 ( .B(fifo_array[771]), .A(fifo_array[805]), .S(n4619), .Y(n4224) );
  MUX2X1 U4569 ( .B(fifo_array[703]), .A(fifo_array[737]), .S(n4619), .Y(n4223) );
  MUX2X1 U4570 ( .B(fifo_array[635]), .A(fifo_array[669]), .S(n4619), .Y(n4227) );
  MUX2X1 U4571 ( .B(fifo_array[567]), .A(fifo_array[601]), .S(n4619), .Y(n4226) );
  MUX2X1 U4572 ( .B(n4225), .A(n4222), .S(n21), .Y(n4229) );
  MUX2X1 U4573 ( .B(fifo_array[499]), .A(fifo_array[533]), .S(n4620), .Y(n4233) );
  MUX2X1 U4574 ( .B(fifo_array[431]), .A(fifo_array[465]), .S(n4620), .Y(n4232) );
  MUX2X1 U4575 ( .B(fifo_array[363]), .A(fifo_array[397]), .S(n4620), .Y(n4236) );
  MUX2X1 U4576 ( .B(fifo_array[295]), .A(fifo_array[329]), .S(n4620), .Y(n4235) );
  MUX2X1 U4577 ( .B(n4234), .A(n4231), .S(n4654), .Y(n4245) );
  MUX2X1 U4578 ( .B(fifo_array[227]), .A(fifo_array[261]), .S(n4620), .Y(n4239) );
  MUX2X1 U4579 ( .B(fifo_array[159]), .A(fifo_array[193]), .S(n4620), .Y(n4238) );
  MUX2X1 U4580 ( .B(fifo_array[91]), .A(fifo_array[125]), .S(n4620), .Y(n4242)
         );
  MUX2X1 U4581 ( .B(fifo_array[23]), .A(fifo_array[57]), .S(n4620), .Y(n4241)
         );
  MUX2X1 U4582 ( .B(n4240), .A(n4237), .S(n21), .Y(n4244) );
  MUX2X1 U4583 ( .B(n4243), .A(n4228), .S(n23), .Y(n4569) );
  MUX2X1 U4584 ( .B(fifo_array[1044]), .A(fifo_array[1078]), .S(n4620), .Y(
        n4248) );
  MUX2X1 U4585 ( .B(fifo_array[976]), .A(fifo_array[1010]), .S(n4620), .Y(
        n4247) );
  MUX2X1 U4586 ( .B(fifo_array[908]), .A(fifo_array[942]), .S(n4620), .Y(n4251) );
  MUX2X1 U4587 ( .B(fifo_array[840]), .A(fifo_array[874]), .S(n4620), .Y(n4250) );
  MUX2X1 U4588 ( .B(n4249), .A(n4246), .S(n4655), .Y(n4260) );
  MUX2X1 U4589 ( .B(fifo_array[772]), .A(fifo_array[806]), .S(n4621), .Y(n4254) );
  MUX2X1 U4590 ( .B(fifo_array[704]), .A(fifo_array[738]), .S(n4621), .Y(n4253) );
  MUX2X1 U4591 ( .B(fifo_array[636]), .A(fifo_array[670]), .S(n4621), .Y(n4257) );
  MUX2X1 U4592 ( .B(fifo_array[568]), .A(fifo_array[602]), .S(n4621), .Y(n4256) );
  MUX2X1 U4593 ( .B(n4255), .A(n4252), .S(n21), .Y(n4259) );
  MUX2X1 U4594 ( .B(fifo_array[500]), .A(fifo_array[534]), .S(n4621), .Y(n4263) );
  MUX2X1 U4595 ( .B(fifo_array[432]), .A(fifo_array[466]), .S(n4621), .Y(n4262) );
  MUX2X1 U4596 ( .B(fifo_array[364]), .A(fifo_array[398]), .S(n4621), .Y(n4266) );
  MUX2X1 U4597 ( .B(fifo_array[296]), .A(fifo_array[330]), .S(n4621), .Y(n4265) );
  MUX2X1 U4598 ( .B(n4264), .A(n4261), .S(n4655), .Y(n4275) );
  MUX2X1 U4599 ( .B(fifo_array[228]), .A(fifo_array[262]), .S(n4621), .Y(n4269) );
  MUX2X1 U4600 ( .B(fifo_array[160]), .A(fifo_array[194]), .S(n4621), .Y(n4268) );
  MUX2X1 U4601 ( .B(fifo_array[92]), .A(fifo_array[126]), .S(n4621), .Y(n4272)
         );
  MUX2X1 U4602 ( .B(fifo_array[24]), .A(fifo_array[58]), .S(n4621), .Y(n4271)
         );
  MUX2X1 U4603 ( .B(n4270), .A(n4267), .S(n21), .Y(n4274) );
  MUX2X1 U4604 ( .B(n4273), .A(n4258), .S(n23), .Y(n4570) );
  MUX2X1 U4605 ( .B(fifo_array[1045]), .A(fifo_array[1079]), .S(n4622), .Y(
        n4278) );
  MUX2X1 U4606 ( .B(fifo_array[977]), .A(fifo_array[1011]), .S(n4622), .Y(
        n4277) );
  MUX2X1 U4607 ( .B(fifo_array[909]), .A(fifo_array[943]), .S(n4622), .Y(n4281) );
  MUX2X1 U4608 ( .B(fifo_array[841]), .A(fifo_array[875]), .S(n4622), .Y(n4280) );
  MUX2X1 U4609 ( .B(n4279), .A(n4276), .S(n21), .Y(n4290) );
  MUX2X1 U4610 ( .B(fifo_array[773]), .A(fifo_array[807]), .S(n4622), .Y(n4284) );
  MUX2X1 U4611 ( .B(fifo_array[705]), .A(fifo_array[739]), .S(n4622), .Y(n4283) );
  MUX2X1 U4612 ( .B(fifo_array[637]), .A(fifo_array[671]), .S(n4622), .Y(n4287) );
  MUX2X1 U4613 ( .B(fifo_array[569]), .A(fifo_array[603]), .S(n4622), .Y(n4286) );
  MUX2X1 U4614 ( .B(n4285), .A(n4282), .S(n21), .Y(n4289) );
  MUX2X1 U4615 ( .B(fifo_array[501]), .A(fifo_array[535]), .S(n4622), .Y(n4293) );
  MUX2X1 U4616 ( .B(fifo_array[433]), .A(fifo_array[467]), .S(n4622), .Y(n4292) );
  MUX2X1 U4617 ( .B(fifo_array[365]), .A(fifo_array[399]), .S(n4622), .Y(n4296) );
  MUX2X1 U4618 ( .B(fifo_array[297]), .A(fifo_array[331]), .S(n4622), .Y(n4295) );
  MUX2X1 U4619 ( .B(n4294), .A(n4291), .S(n21), .Y(n4305) );
  MUX2X1 U4620 ( .B(fifo_array[229]), .A(fifo_array[263]), .S(n4623), .Y(n4299) );
  MUX2X1 U4621 ( .B(fifo_array[161]), .A(fifo_array[195]), .S(n4623), .Y(n4298) );
  MUX2X1 U4622 ( .B(fifo_array[93]), .A(fifo_array[127]), .S(n4623), .Y(n4302)
         );
  MUX2X1 U4623 ( .B(fifo_array[25]), .A(fifo_array[59]), .S(n4623), .Y(n4301)
         );
  MUX2X1 U4624 ( .B(n4300), .A(n4297), .S(n21), .Y(n4304) );
  MUX2X1 U4625 ( .B(n4303), .A(n4288), .S(n23), .Y(n4571) );
  MUX2X1 U4626 ( .B(fifo_array[1046]), .A(fifo_array[1080]), .S(n4623), .Y(
        n4308) );
  MUX2X1 U4627 ( .B(fifo_array[978]), .A(fifo_array[1012]), .S(n4623), .Y(
        n4307) );
  MUX2X1 U4628 ( .B(fifo_array[910]), .A(fifo_array[944]), .S(n4623), .Y(n4311) );
  MUX2X1 U4629 ( .B(fifo_array[842]), .A(fifo_array[876]), .S(n4623), .Y(n4310) );
  MUX2X1 U4630 ( .B(n4309), .A(n4306), .S(n21), .Y(n4320) );
  MUX2X1 U4631 ( .B(fifo_array[774]), .A(fifo_array[808]), .S(n4623), .Y(n4314) );
  MUX2X1 U4632 ( .B(fifo_array[706]), .A(fifo_array[740]), .S(n4623), .Y(n4313) );
  MUX2X1 U4633 ( .B(fifo_array[638]), .A(fifo_array[672]), .S(n4623), .Y(n4317) );
  MUX2X1 U4634 ( .B(fifo_array[570]), .A(fifo_array[604]), .S(n4623), .Y(n4316) );
  MUX2X1 U4635 ( .B(n4315), .A(n4312), .S(n21), .Y(n4319) );
  MUX2X1 U4636 ( .B(fifo_array[502]), .A(fifo_array[536]), .S(n4624), .Y(n4323) );
  MUX2X1 U4637 ( .B(fifo_array[434]), .A(fifo_array[468]), .S(n4624), .Y(n4322) );
  MUX2X1 U4638 ( .B(fifo_array[366]), .A(fifo_array[400]), .S(n4624), .Y(n4326) );
  MUX2X1 U4639 ( .B(fifo_array[298]), .A(fifo_array[332]), .S(n4624), .Y(n4325) );
  MUX2X1 U4640 ( .B(n4324), .A(n4321), .S(n21), .Y(n4335) );
  MUX2X1 U4641 ( .B(fifo_array[230]), .A(fifo_array[264]), .S(n4624), .Y(n4329) );
  MUX2X1 U4642 ( .B(fifo_array[162]), .A(fifo_array[196]), .S(n4624), .Y(n4328) );
  MUX2X1 U4643 ( .B(fifo_array[94]), .A(fifo_array[128]), .S(n4624), .Y(n4332)
         );
  MUX2X1 U4644 ( .B(fifo_array[26]), .A(fifo_array[60]), .S(n4624), .Y(n4331)
         );
  MUX2X1 U4645 ( .B(n4330), .A(n4327), .S(n21), .Y(n4334) );
  MUX2X1 U4646 ( .B(n4333), .A(n4318), .S(n23), .Y(n4572) );
  MUX2X1 U4647 ( .B(fifo_array[1047]), .A(fifo_array[1081]), .S(n4624), .Y(
        n4338) );
  MUX2X1 U4648 ( .B(fifo_array[979]), .A(fifo_array[1013]), .S(n4624), .Y(
        n4337) );
  MUX2X1 U4649 ( .B(fifo_array[911]), .A(fifo_array[945]), .S(n4624), .Y(n4341) );
  MUX2X1 U4650 ( .B(fifo_array[843]), .A(fifo_array[877]), .S(n4624), .Y(n4340) );
  MUX2X1 U4651 ( .B(n4339), .A(n4336), .S(n21), .Y(n4350) );
  MUX2X1 U4652 ( .B(fifo_array[775]), .A(fifo_array[809]), .S(n4625), .Y(n4344) );
  MUX2X1 U4653 ( .B(fifo_array[707]), .A(fifo_array[741]), .S(n4625), .Y(n4343) );
  MUX2X1 U4654 ( .B(fifo_array[639]), .A(fifo_array[673]), .S(n4625), .Y(n4347) );
  MUX2X1 U4655 ( .B(fifo_array[571]), .A(fifo_array[605]), .S(n4625), .Y(n4346) );
  MUX2X1 U4656 ( .B(n4345), .A(n4342), .S(n21), .Y(n4349) );
  MUX2X1 U4657 ( .B(fifo_array[503]), .A(fifo_array[537]), .S(n4625), .Y(n4353) );
  MUX2X1 U4658 ( .B(fifo_array[435]), .A(fifo_array[469]), .S(n4625), .Y(n4352) );
  MUX2X1 U4659 ( .B(fifo_array[367]), .A(fifo_array[401]), .S(n4625), .Y(n4356) );
  MUX2X1 U4660 ( .B(fifo_array[299]), .A(fifo_array[333]), .S(n4625), .Y(n4355) );
  MUX2X1 U4661 ( .B(n4354), .A(n4351), .S(n21), .Y(n4365) );
  MUX2X1 U4662 ( .B(fifo_array[231]), .A(fifo_array[265]), .S(n4625), .Y(n4359) );
  MUX2X1 U4663 ( .B(fifo_array[163]), .A(fifo_array[197]), .S(n4625), .Y(n4358) );
  MUX2X1 U4664 ( .B(fifo_array[95]), .A(fifo_array[129]), .S(n4625), .Y(n4362)
         );
  MUX2X1 U4665 ( .B(fifo_array[27]), .A(fifo_array[61]), .S(n4625), .Y(n4361)
         );
  MUX2X1 U4666 ( .B(n4360), .A(n4357), .S(n21), .Y(n4364) );
  MUX2X1 U4667 ( .B(n4363), .A(n4348), .S(n23), .Y(n4573) );
  MUX2X1 U4668 ( .B(fifo_array[1048]), .A(fifo_array[1082]), .S(n4626), .Y(
        n4368) );
  MUX2X1 U4669 ( .B(fifo_array[980]), .A(fifo_array[1014]), .S(n4626), .Y(
        n4367) );
  MUX2X1 U4670 ( .B(fifo_array[912]), .A(fifo_array[946]), .S(n4626), .Y(n4371) );
  MUX2X1 U4671 ( .B(fifo_array[844]), .A(fifo_array[878]), .S(n4626), .Y(n4370) );
  MUX2X1 U4672 ( .B(n4369), .A(n4366), .S(n21), .Y(n4380) );
  MUX2X1 U4673 ( .B(fifo_array[776]), .A(fifo_array[810]), .S(n4626), .Y(n4374) );
  MUX2X1 U4674 ( .B(fifo_array[708]), .A(fifo_array[742]), .S(n4626), .Y(n4373) );
  MUX2X1 U4675 ( .B(fifo_array[640]), .A(fifo_array[674]), .S(n4626), .Y(n4377) );
  MUX2X1 U4676 ( .B(fifo_array[572]), .A(fifo_array[606]), .S(n4626), .Y(n4376) );
  MUX2X1 U4677 ( .B(n4375), .A(n4372), .S(n21), .Y(n4379) );
  MUX2X1 U4678 ( .B(fifo_array[504]), .A(fifo_array[538]), .S(n4626), .Y(n4383) );
  MUX2X1 U4679 ( .B(fifo_array[436]), .A(fifo_array[470]), .S(n4626), .Y(n4382) );
  MUX2X1 U4680 ( .B(fifo_array[368]), .A(fifo_array[402]), .S(n4626), .Y(n4386) );
  MUX2X1 U4681 ( .B(fifo_array[300]), .A(fifo_array[334]), .S(n4626), .Y(n4385) );
  MUX2X1 U4682 ( .B(n4384), .A(n4381), .S(n21), .Y(n4395) );
  MUX2X1 U4683 ( .B(fifo_array[232]), .A(fifo_array[266]), .S(n4627), .Y(n4389) );
  MUX2X1 U4684 ( .B(fifo_array[164]), .A(fifo_array[198]), .S(n4627), .Y(n4388) );
  MUX2X1 U4685 ( .B(fifo_array[96]), .A(fifo_array[130]), .S(n4627), .Y(n4392)
         );
  MUX2X1 U4686 ( .B(fifo_array[28]), .A(fifo_array[62]), .S(n4627), .Y(n4391)
         );
  MUX2X1 U4687 ( .B(n4390), .A(n4387), .S(n21), .Y(n4394) );
  MUX2X1 U4688 ( .B(n4393), .A(n4378), .S(n23), .Y(n4574) );
  MUX2X1 U4689 ( .B(fifo_array[1049]), .A(fifo_array[1083]), .S(n4627), .Y(
        n4398) );
  MUX2X1 U4690 ( .B(fifo_array[981]), .A(fifo_array[1015]), .S(n4627), .Y(
        n4397) );
  MUX2X1 U4691 ( .B(fifo_array[913]), .A(fifo_array[947]), .S(n4627), .Y(n4401) );
  MUX2X1 U4692 ( .B(fifo_array[845]), .A(fifo_array[879]), .S(n4627), .Y(n4400) );
  MUX2X1 U4693 ( .B(n4399), .A(n4396), .S(n21), .Y(n4410) );
  MUX2X1 U4694 ( .B(fifo_array[777]), .A(fifo_array[811]), .S(n4627), .Y(n4404) );
  MUX2X1 U4695 ( .B(fifo_array[709]), .A(fifo_array[743]), .S(n4627), .Y(n4403) );
  MUX2X1 U4696 ( .B(fifo_array[641]), .A(fifo_array[675]), .S(n4627), .Y(n4407) );
  MUX2X1 U4697 ( .B(fifo_array[573]), .A(fifo_array[607]), .S(n4627), .Y(n4406) );
  MUX2X1 U4698 ( .B(n4405), .A(n4402), .S(n21), .Y(n4409) );
  MUX2X1 U4699 ( .B(fifo_array[505]), .A(fifo_array[539]), .S(n4628), .Y(n4413) );
  MUX2X1 U4700 ( .B(fifo_array[437]), .A(fifo_array[471]), .S(n4628), .Y(n4412) );
  MUX2X1 U4701 ( .B(fifo_array[369]), .A(fifo_array[403]), .S(n4628), .Y(n4416) );
  MUX2X1 U4702 ( .B(fifo_array[301]), .A(fifo_array[335]), .S(n4628), .Y(n4415) );
  MUX2X1 U4703 ( .B(n4414), .A(n4411), .S(n21), .Y(n4425) );
  MUX2X1 U4704 ( .B(fifo_array[233]), .A(fifo_array[267]), .S(n4628), .Y(n4419) );
  MUX2X1 U4705 ( .B(fifo_array[165]), .A(fifo_array[199]), .S(n4628), .Y(n4418) );
  MUX2X1 U4706 ( .B(fifo_array[97]), .A(fifo_array[131]), .S(n4628), .Y(n4422)
         );
  MUX2X1 U4707 ( .B(fifo_array[29]), .A(fifo_array[63]), .S(n4628), .Y(n4421)
         );
  MUX2X1 U4708 ( .B(n4420), .A(n4417), .S(n21), .Y(n4424) );
  MUX2X1 U4709 ( .B(n4423), .A(n4408), .S(n23), .Y(n4575) );
  MUX2X1 U4710 ( .B(fifo_array[1050]), .A(fifo_array[1084]), .S(n4628), .Y(
        n4428) );
  MUX2X1 U4711 ( .B(fifo_array[982]), .A(fifo_array[1016]), .S(n4628), .Y(
        n4427) );
  MUX2X1 U4712 ( .B(fifo_array[914]), .A(fifo_array[948]), .S(n4628), .Y(n4431) );
  MUX2X1 U4713 ( .B(fifo_array[846]), .A(fifo_array[880]), .S(n4628), .Y(n4430) );
  MUX2X1 U4714 ( .B(n4429), .A(n4426), .S(n21), .Y(n4440) );
  MUX2X1 U4715 ( .B(fifo_array[778]), .A(fifo_array[812]), .S(n4629), .Y(n4434) );
  MUX2X1 U4716 ( .B(fifo_array[710]), .A(fifo_array[744]), .S(n4629), .Y(n4433) );
  MUX2X1 U4717 ( .B(fifo_array[642]), .A(fifo_array[676]), .S(n4629), .Y(n4437) );
  MUX2X1 U4718 ( .B(fifo_array[574]), .A(fifo_array[608]), .S(n4629), .Y(n4436) );
  MUX2X1 U4719 ( .B(n4435), .A(n4432), .S(n21), .Y(n4439) );
  MUX2X1 U4720 ( .B(fifo_array[506]), .A(fifo_array[540]), .S(n4629), .Y(n4443) );
  MUX2X1 U4721 ( .B(fifo_array[438]), .A(fifo_array[472]), .S(n4629), .Y(n4442) );
  MUX2X1 U4722 ( .B(fifo_array[370]), .A(fifo_array[404]), .S(n4629), .Y(n4446) );
  MUX2X1 U4723 ( .B(fifo_array[302]), .A(fifo_array[336]), .S(n4629), .Y(n4445) );
  MUX2X1 U4724 ( .B(n4444), .A(n4441), .S(n21), .Y(n4455) );
  MUX2X1 U4725 ( .B(fifo_array[234]), .A(fifo_array[268]), .S(n4629), .Y(n4449) );
  MUX2X1 U4726 ( .B(fifo_array[166]), .A(fifo_array[200]), .S(n4629), .Y(n4448) );
  MUX2X1 U4727 ( .B(fifo_array[98]), .A(fifo_array[132]), .S(n4629), .Y(n4452)
         );
  MUX2X1 U4728 ( .B(fifo_array[30]), .A(fifo_array[64]), .S(n4629), .Y(n4451)
         );
  MUX2X1 U4729 ( .B(n4450), .A(n4447), .S(n21), .Y(n4454) );
  MUX2X1 U4730 ( .B(n4453), .A(n4438), .S(n23), .Y(n4576) );
  MUX2X1 U4731 ( .B(fifo_array[1051]), .A(fifo_array[1085]), .S(n4630), .Y(
        n4458) );
  MUX2X1 U4732 ( .B(fifo_array[983]), .A(fifo_array[1017]), .S(n4630), .Y(
        n4457) );
  MUX2X1 U4733 ( .B(fifo_array[915]), .A(fifo_array[949]), .S(n4630), .Y(n4461) );
  MUX2X1 U4734 ( .B(fifo_array[847]), .A(fifo_array[881]), .S(n4630), .Y(n4460) );
  MUX2X1 U4735 ( .B(n4459), .A(n4456), .S(n21), .Y(n4470) );
  MUX2X1 U4736 ( .B(fifo_array[779]), .A(fifo_array[813]), .S(n4630), .Y(n4464) );
  MUX2X1 U4737 ( .B(fifo_array[711]), .A(fifo_array[745]), .S(n4630), .Y(n4463) );
  MUX2X1 U4738 ( .B(fifo_array[643]), .A(fifo_array[677]), .S(n4630), .Y(n4467) );
  MUX2X1 U4739 ( .B(fifo_array[575]), .A(fifo_array[609]), .S(n4630), .Y(n4466) );
  MUX2X1 U4740 ( .B(n4465), .A(n4462), .S(n21), .Y(n4469) );
  MUX2X1 U4741 ( .B(fifo_array[507]), .A(fifo_array[541]), .S(n4630), .Y(n4473) );
  MUX2X1 U4742 ( .B(fifo_array[439]), .A(fifo_array[473]), .S(n4630), .Y(n4472) );
  MUX2X1 U4743 ( .B(fifo_array[371]), .A(fifo_array[405]), .S(n4630), .Y(n4476) );
  MUX2X1 U4744 ( .B(fifo_array[303]), .A(fifo_array[337]), .S(n4630), .Y(n4475) );
  MUX2X1 U4745 ( .B(n4474), .A(n4471), .S(n21), .Y(n4485) );
  MUX2X1 U4746 ( .B(fifo_array[235]), .A(fifo_array[269]), .S(n4631), .Y(n4479) );
  MUX2X1 U4747 ( .B(fifo_array[167]), .A(fifo_array[201]), .S(n4631), .Y(n4478) );
  MUX2X1 U4748 ( .B(fifo_array[99]), .A(fifo_array[133]), .S(n4631), .Y(n4482)
         );
  MUX2X1 U4749 ( .B(fifo_array[31]), .A(fifo_array[65]), .S(n4631), .Y(n4481)
         );
  MUX2X1 U4750 ( .B(n4480), .A(n4477), .S(n21), .Y(n4484) );
  MUX2X1 U4751 ( .B(n4483), .A(n4468), .S(n23), .Y(n4577) );
  MUX2X1 U4752 ( .B(fifo_array[1052]), .A(fifo_array[1086]), .S(n4631), .Y(
        n4488) );
  MUX2X1 U4753 ( .B(fifo_array[984]), .A(fifo_array[1018]), .S(n4631), .Y(
        n4487) );
  MUX2X1 U4754 ( .B(fifo_array[916]), .A(fifo_array[950]), .S(n4631), .Y(n4491) );
  MUX2X1 U4755 ( .B(fifo_array[848]), .A(fifo_array[882]), .S(n4631), .Y(n4490) );
  MUX2X1 U4756 ( .B(n4489), .A(n4486), .S(n21), .Y(n4500) );
  MUX2X1 U4757 ( .B(fifo_array[780]), .A(fifo_array[814]), .S(n4631), .Y(n4494) );
  MUX2X1 U4758 ( .B(fifo_array[712]), .A(fifo_array[746]), .S(n4631), .Y(n4493) );
  MUX2X1 U4759 ( .B(fifo_array[644]), .A(fifo_array[678]), .S(n4631), .Y(n4497) );
  MUX2X1 U4760 ( .B(fifo_array[576]), .A(fifo_array[610]), .S(n4631), .Y(n4496) );
  MUX2X1 U4761 ( .B(n4495), .A(n4492), .S(n21), .Y(n4499) );
  MUX2X1 U4762 ( .B(fifo_array[508]), .A(fifo_array[542]), .S(n4632), .Y(n4503) );
  MUX2X1 U4763 ( .B(fifo_array[440]), .A(fifo_array[474]), .S(n4632), .Y(n4502) );
  MUX2X1 U4764 ( .B(fifo_array[372]), .A(fifo_array[406]), .S(n4632), .Y(n4506) );
  MUX2X1 U4765 ( .B(fifo_array[304]), .A(fifo_array[338]), .S(n4632), .Y(n4505) );
  MUX2X1 U4766 ( .B(n4504), .A(n4501), .S(n21), .Y(n4515) );
  MUX2X1 U4767 ( .B(fifo_array[236]), .A(fifo_array[270]), .S(n4632), .Y(n4509) );
  MUX2X1 U4768 ( .B(fifo_array[168]), .A(fifo_array[202]), .S(n4632), .Y(n4508) );
  MUX2X1 U4769 ( .B(fifo_array[100]), .A(fifo_array[134]), .S(n4632), .Y(n4512) );
  MUX2X1 U4770 ( .B(fifo_array[32]), .A(fifo_array[66]), .S(n4632), .Y(n4511)
         );
  MUX2X1 U4771 ( .B(n4510), .A(n4507), .S(n21), .Y(n4514) );
  MUX2X1 U4772 ( .B(n4513), .A(n4498), .S(n23), .Y(n4578) );
  MUX2X1 U4773 ( .B(fifo_array[1053]), .A(fifo_array[1087]), .S(n4632), .Y(
        n4518) );
  MUX2X1 U4774 ( .B(fifo_array[985]), .A(fifo_array[1019]), .S(n4632), .Y(
        n4517) );
  MUX2X1 U4775 ( .B(fifo_array[917]), .A(fifo_array[951]), .S(n4632), .Y(n4521) );
  MUX2X1 U4776 ( .B(fifo_array[849]), .A(fifo_array[883]), .S(n4632), .Y(n4520) );
  MUX2X1 U4777 ( .B(n4519), .A(n4516), .S(n21), .Y(n4530) );
  MUX2X1 U4778 ( .B(fifo_array[781]), .A(fifo_array[815]), .S(n4633), .Y(n4524) );
  MUX2X1 U4779 ( .B(fifo_array[713]), .A(fifo_array[747]), .S(n4633), .Y(n4523) );
  MUX2X1 U4780 ( .B(fifo_array[645]), .A(fifo_array[679]), .S(n4633), .Y(n4527) );
  MUX2X1 U4781 ( .B(fifo_array[577]), .A(fifo_array[611]), .S(n4633), .Y(n4526) );
  MUX2X1 U4782 ( .B(n4525), .A(n4522), .S(n21), .Y(n4529) );
  MUX2X1 U4783 ( .B(fifo_array[509]), .A(fifo_array[543]), .S(n4633), .Y(n4533) );
  MUX2X1 U4784 ( .B(fifo_array[441]), .A(fifo_array[475]), .S(n4633), .Y(n4532) );
  MUX2X1 U4785 ( .B(fifo_array[373]), .A(fifo_array[407]), .S(n4633), .Y(n4536) );
  MUX2X1 U4786 ( .B(fifo_array[305]), .A(fifo_array[339]), .S(n4633), .Y(n4535) );
  MUX2X1 U4787 ( .B(n4534), .A(n4531), .S(n21), .Y(n4545) );
  MUX2X1 U4788 ( .B(fifo_array[237]), .A(fifo_array[271]), .S(n4633), .Y(n4539) );
  MUX2X1 U4789 ( .B(fifo_array[169]), .A(fifo_array[203]), .S(n4633), .Y(n4538) );
  MUX2X1 U4790 ( .B(fifo_array[101]), .A(fifo_array[135]), .S(n4633), .Y(n4542) );
  MUX2X1 U4791 ( .B(fifo_array[33]), .A(fifo_array[67]), .S(n4633), .Y(n4541)
         );
  MUX2X1 U4792 ( .B(n4540), .A(n4537), .S(n21), .Y(n4544) );
  MUX2X1 U4793 ( .B(n4543), .A(n4528), .S(n23), .Y(n4579) );
  XOR2X1 U4794 ( .A(r307_carry[4]), .B(wr_ptr[4]), .Y(n71) );
  XOR2X1 U4795 ( .A(r308_carry[4]), .B(n23), .Y(n76) );
  XOR2X1 U4796 ( .A(add_45_carry[5]), .B(fillcount[5]), .Y(n88) );
  OAI21X1 U4797 ( .A(n95), .B(n4814), .C(n3521), .Y(n96) );
  OAI21X1 U4798 ( .A(n4759), .B(n4764), .C(n3455), .Y(n97) );
  OAI21X1 U4799 ( .A(n4760), .B(n4763), .C(n3522), .Y(n98) );
  XNOR2X1 U4800 ( .A(fillcount[4]), .B(n3522), .Y(n99) );
  XNOR2X1 U4801 ( .A(fillcount[5]), .B(n4762), .Y(n100) );
endmodule


module FIFO_DEPTH_P25_WIDTH42 ( clk, reset, data_in, put, get, data_out, empty, 
        full, fillcount );
  input [41:0] data_in;
  output [41:0] data_out;
  output [5:0] fillcount;
  input clk, reset, put, get;
  output empty, full;
  wire   n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n76, n77, n78, n79, n81, n82, n83, n84, n92,
         n93, n94, n95, n96, n103, n104, n105, n106, n107, n108, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n80, n85, n86, n87, n88, n89,
         n90, n91, n97, n98, n99, n100, n101, n102, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n1585,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904;
  wire   [4:0] wr_ptr;
  wire   [1343:0] fifo_array;
  wire   [5:2] add_45_carry;
  wire   [4:2] r308_carry;
  wire   [4:2] r307_carry;

  DFFPOSX1 full_reg ( .D(n3012), .CLK(clk), .Q(full) );
  DFFPOSX1 fillcount_reg_5_ ( .D(n3011), .CLK(clk), .Q(fillcount[5]) );
  DFFPOSX1 empty_reg ( .D(n3010), .CLK(clk), .Q(empty) );
  DFFPOSX1 wr_ptr_reg_0_ ( .D(n2999), .CLK(clk), .Q(wr_ptr[0]) );
  DFFPOSX1 wr_ptr_reg_1_ ( .D(n2998), .CLK(clk), .Q(wr_ptr[1]) );
  DFFPOSX1 wr_ptr_reg_2_ ( .D(n2997), .CLK(clk), .Q(wr_ptr[2]) );
  DFFPOSX1 wr_ptr_reg_3_ ( .D(n2996), .CLK(clk), .Q(wr_ptr[3]) );
  DFFPOSX1 wr_ptr_reg_4_ ( .D(n2995), .CLK(clk), .Q(wr_ptr[4]) );
  DFFPOSX1 data_out_reg_0_ ( .D(n5852), .CLK(clk), .Q(data_out[0]) );
  DFFPOSX1 data_out_reg_1_ ( .D(n5853), .CLK(clk), .Q(data_out[1]) );
  DFFPOSX1 data_out_reg_2_ ( .D(n5854), .CLK(clk), .Q(data_out[2]) );
  DFFPOSX1 data_out_reg_3_ ( .D(n5855), .CLK(clk), .Q(data_out[3]) );
  DFFPOSX1 data_out_reg_4_ ( .D(n5856), .CLK(clk), .Q(data_out[4]) );
  DFFPOSX1 data_out_reg_5_ ( .D(n5857), .CLK(clk), .Q(data_out[5]) );
  DFFPOSX1 data_out_reg_6_ ( .D(n5858), .CLK(clk), .Q(data_out[6]) );
  DFFPOSX1 data_out_reg_7_ ( .D(n5859), .CLK(clk), .Q(data_out[7]) );
  DFFPOSX1 data_out_reg_8_ ( .D(n5860), .CLK(clk), .Q(data_out[8]) );
  DFFPOSX1 data_out_reg_9_ ( .D(n5861), .CLK(clk), .Q(data_out[9]) );
  DFFPOSX1 data_out_reg_10_ ( .D(n5862), .CLK(clk), .Q(data_out[10]) );
  DFFPOSX1 data_out_reg_11_ ( .D(n5863), .CLK(clk), .Q(data_out[11]) );
  DFFPOSX1 data_out_reg_12_ ( .D(n5864), .CLK(clk), .Q(data_out[12]) );
  DFFPOSX1 data_out_reg_13_ ( .D(n5865), .CLK(clk), .Q(data_out[13]) );
  DFFPOSX1 data_out_reg_14_ ( .D(n5866), .CLK(clk), .Q(data_out[14]) );
  DFFPOSX1 data_out_reg_15_ ( .D(n5867), .CLK(clk), .Q(data_out[15]) );
  DFFPOSX1 data_out_reg_16_ ( .D(n5868), .CLK(clk), .Q(data_out[16]) );
  DFFPOSX1 data_out_reg_17_ ( .D(n5869), .CLK(clk), .Q(data_out[17]) );
  DFFPOSX1 data_out_reg_18_ ( .D(n5870), .CLK(clk), .Q(data_out[18]) );
  DFFPOSX1 data_out_reg_19_ ( .D(n5871), .CLK(clk), .Q(data_out[19]) );
  DFFPOSX1 data_out_reg_20_ ( .D(n5872), .CLK(clk), .Q(data_out[20]) );
  DFFPOSX1 data_out_reg_21_ ( .D(n5873), .CLK(clk), .Q(data_out[21]) );
  DFFPOSX1 data_out_reg_22_ ( .D(n5874), .CLK(clk), .Q(data_out[22]) );
  DFFPOSX1 data_out_reg_23_ ( .D(n5875), .CLK(clk), .Q(data_out[23]) );
  DFFPOSX1 data_out_reg_24_ ( .D(n5876), .CLK(clk), .Q(data_out[24]) );
  DFFPOSX1 data_out_reg_25_ ( .D(n5877), .CLK(clk), .Q(data_out[25]) );
  DFFPOSX1 data_out_reg_26_ ( .D(n5878), .CLK(clk), .Q(data_out[26]) );
  DFFPOSX1 data_out_reg_27_ ( .D(n5879), .CLK(clk), .Q(data_out[27]) );
  DFFPOSX1 data_out_reg_28_ ( .D(n5880), .CLK(clk), .Q(data_out[28]) );
  DFFPOSX1 data_out_reg_29_ ( .D(n5881), .CLK(clk), .Q(data_out[29]) );
  DFFPOSX1 data_out_reg_30_ ( .D(n5882), .CLK(clk), .Q(data_out[30]) );
  DFFPOSX1 data_out_reg_31_ ( .D(n5883), .CLK(clk), .Q(data_out[31]) );
  DFFPOSX1 data_out_reg_32_ ( .D(n5884), .CLK(clk), .Q(data_out[32]) );
  DFFPOSX1 data_out_reg_33_ ( .D(n5885), .CLK(clk), .Q(data_out[33]) );
  DFFPOSX1 data_out_reg_34_ ( .D(n5886), .CLK(clk), .Q(data_out[34]) );
  DFFPOSX1 data_out_reg_35_ ( .D(n5887), .CLK(clk), .Q(data_out[35]) );
  DFFPOSX1 data_out_reg_36_ ( .D(n5888), .CLK(clk), .Q(data_out[36]) );
  DFFPOSX1 data_out_reg_37_ ( .D(n5889), .CLK(clk), .Q(data_out[37]) );
  DFFPOSX1 data_out_reg_38_ ( .D(n5890), .CLK(clk), .Q(data_out[38]) );
  DFFPOSX1 data_out_reg_39_ ( .D(n5891), .CLK(clk), .Q(data_out[39]) );
  DFFPOSX1 data_out_reg_40_ ( .D(n5892), .CLK(clk), .Q(data_out[40]) );
  DFFPOSX1 data_out_reg_41_ ( .D(n5893), .CLK(clk), .Q(data_out[41]) );
  DFFPOSX1 rd_ptr_reg_0_ ( .D(n3009), .CLK(clk), .Q(n19) );
  DFFPOSX1 rd_ptr_reg_1_ ( .D(n3008), .CLK(clk), .Q(n20) );
  DFFPOSX1 rd_ptr_reg_2_ ( .D(n3007), .CLK(clk), .Q(n21) );
  DFFPOSX1 rd_ptr_reg_3_ ( .D(n3006), .CLK(clk), .Q(n22) );
  DFFPOSX1 rd_ptr_reg_4_ ( .D(n3005), .CLK(clk), .Q(n23) );
  DFFPOSX1 fillcount_reg_0_ ( .D(n3004), .CLK(clk), .Q(fillcount[0]) );
  DFFPOSX1 fillcount_reg_4_ ( .D(n3000), .CLK(clk), .Q(fillcount[4]) );
  DFFPOSX1 fillcount_reg_1_ ( .D(n3003), .CLK(clk), .Q(fillcount[1]) );
  DFFPOSX1 fillcount_reg_2_ ( .D(n3002), .CLK(clk), .Q(fillcount[2]) );
  DFFPOSX1 fillcount_reg_3_ ( .D(n3001), .CLK(clk), .Q(fillcount[3]) );
  DFFPOSX1 fifo_array_reg_31__41_ ( .D(n2994), .CLK(clk), .Q(fifo_array[1343])
         );
  DFFPOSX1 fifo_array_reg_31__40_ ( .D(n2993), .CLK(clk), .Q(fifo_array[1342])
         );
  DFFPOSX1 fifo_array_reg_31__39_ ( .D(n2992), .CLK(clk), .Q(fifo_array[1341])
         );
  DFFPOSX1 fifo_array_reg_31__38_ ( .D(n2991), .CLK(clk), .Q(fifo_array[1340])
         );
  DFFPOSX1 fifo_array_reg_31__37_ ( .D(n2990), .CLK(clk), .Q(fifo_array[1339])
         );
  DFFPOSX1 fifo_array_reg_31__36_ ( .D(n2989), .CLK(clk), .Q(fifo_array[1338])
         );
  DFFPOSX1 fifo_array_reg_31__35_ ( .D(n2988), .CLK(clk), .Q(fifo_array[1337])
         );
  DFFPOSX1 fifo_array_reg_31__34_ ( .D(n2987), .CLK(clk), .Q(fifo_array[1336])
         );
  DFFPOSX1 fifo_array_reg_31__33_ ( .D(n2986), .CLK(clk), .Q(fifo_array[1335])
         );
  DFFPOSX1 fifo_array_reg_31__32_ ( .D(n2985), .CLK(clk), .Q(fifo_array[1334])
         );
  DFFPOSX1 fifo_array_reg_31__31_ ( .D(n2984), .CLK(clk), .Q(fifo_array[1333])
         );
  DFFPOSX1 fifo_array_reg_31__30_ ( .D(n2983), .CLK(clk), .Q(fifo_array[1332])
         );
  DFFPOSX1 fifo_array_reg_31__29_ ( .D(n2982), .CLK(clk), .Q(fifo_array[1331])
         );
  DFFPOSX1 fifo_array_reg_31__28_ ( .D(n2981), .CLK(clk), .Q(fifo_array[1330])
         );
  DFFPOSX1 fifo_array_reg_31__27_ ( .D(n2980), .CLK(clk), .Q(fifo_array[1329])
         );
  DFFPOSX1 fifo_array_reg_31__26_ ( .D(n2979), .CLK(clk), .Q(fifo_array[1328])
         );
  DFFPOSX1 fifo_array_reg_31__25_ ( .D(n2978), .CLK(clk), .Q(fifo_array[1327])
         );
  DFFPOSX1 fifo_array_reg_31__24_ ( .D(n2977), .CLK(clk), .Q(fifo_array[1326])
         );
  DFFPOSX1 fifo_array_reg_31__23_ ( .D(n2976), .CLK(clk), .Q(fifo_array[1325])
         );
  DFFPOSX1 fifo_array_reg_31__22_ ( .D(n2975), .CLK(clk), .Q(fifo_array[1324])
         );
  DFFPOSX1 fifo_array_reg_31__21_ ( .D(n2974), .CLK(clk), .Q(fifo_array[1323])
         );
  DFFPOSX1 fifo_array_reg_31__20_ ( .D(n2973), .CLK(clk), .Q(fifo_array[1322])
         );
  DFFPOSX1 fifo_array_reg_31__19_ ( .D(n2972), .CLK(clk), .Q(fifo_array[1321])
         );
  DFFPOSX1 fifo_array_reg_31__18_ ( .D(n2971), .CLK(clk), .Q(fifo_array[1320])
         );
  DFFPOSX1 fifo_array_reg_31__17_ ( .D(n2970), .CLK(clk), .Q(fifo_array[1319])
         );
  DFFPOSX1 fifo_array_reg_31__16_ ( .D(n2969), .CLK(clk), .Q(fifo_array[1318])
         );
  DFFPOSX1 fifo_array_reg_31__15_ ( .D(n2968), .CLK(clk), .Q(fifo_array[1317])
         );
  DFFPOSX1 fifo_array_reg_31__14_ ( .D(n2967), .CLK(clk), .Q(fifo_array[1316])
         );
  DFFPOSX1 fifo_array_reg_31__13_ ( .D(n2966), .CLK(clk), .Q(fifo_array[1315])
         );
  DFFPOSX1 fifo_array_reg_31__12_ ( .D(n2965), .CLK(clk), .Q(fifo_array[1314])
         );
  DFFPOSX1 fifo_array_reg_31__11_ ( .D(n2964), .CLK(clk), .Q(fifo_array[1313])
         );
  DFFPOSX1 fifo_array_reg_31__10_ ( .D(n2963), .CLK(clk), .Q(fifo_array[1312])
         );
  DFFPOSX1 fifo_array_reg_31__9_ ( .D(n2962), .CLK(clk), .Q(fifo_array[1311])
         );
  DFFPOSX1 fifo_array_reg_31__8_ ( .D(n2961), .CLK(clk), .Q(fifo_array[1310])
         );
  DFFPOSX1 fifo_array_reg_31__7_ ( .D(n2960), .CLK(clk), .Q(fifo_array[1309])
         );
  DFFPOSX1 fifo_array_reg_31__6_ ( .D(n2959), .CLK(clk), .Q(fifo_array[1308])
         );
  DFFPOSX1 fifo_array_reg_31__5_ ( .D(n2958), .CLK(clk), .Q(fifo_array[1307])
         );
  DFFPOSX1 fifo_array_reg_31__4_ ( .D(n2957), .CLK(clk), .Q(fifo_array[1306])
         );
  DFFPOSX1 fifo_array_reg_31__3_ ( .D(n2956), .CLK(clk), .Q(fifo_array[1305])
         );
  DFFPOSX1 fifo_array_reg_31__2_ ( .D(n2955), .CLK(clk), .Q(fifo_array[1304])
         );
  DFFPOSX1 fifo_array_reg_31__1_ ( .D(n2954), .CLK(clk), .Q(fifo_array[1303])
         );
  DFFPOSX1 fifo_array_reg_31__0_ ( .D(n2953), .CLK(clk), .Q(fifo_array[1302])
         );
  DFFPOSX1 fifo_array_reg_30__41_ ( .D(n2952), .CLK(clk), .Q(fifo_array[1301])
         );
  DFFPOSX1 fifo_array_reg_30__40_ ( .D(n2951), .CLK(clk), .Q(fifo_array[1300])
         );
  DFFPOSX1 fifo_array_reg_30__39_ ( .D(n2950), .CLK(clk), .Q(fifo_array[1299])
         );
  DFFPOSX1 fifo_array_reg_30__38_ ( .D(n2949), .CLK(clk), .Q(fifo_array[1298])
         );
  DFFPOSX1 fifo_array_reg_30__37_ ( .D(n2948), .CLK(clk), .Q(fifo_array[1297])
         );
  DFFPOSX1 fifo_array_reg_30__36_ ( .D(n2947), .CLK(clk), .Q(fifo_array[1296])
         );
  DFFPOSX1 fifo_array_reg_30__35_ ( .D(n2946), .CLK(clk), .Q(fifo_array[1295])
         );
  DFFPOSX1 fifo_array_reg_30__34_ ( .D(n2945), .CLK(clk), .Q(fifo_array[1294])
         );
  DFFPOSX1 fifo_array_reg_30__33_ ( .D(n2944), .CLK(clk), .Q(fifo_array[1293])
         );
  DFFPOSX1 fifo_array_reg_30__32_ ( .D(n2943), .CLK(clk), .Q(fifo_array[1292])
         );
  DFFPOSX1 fifo_array_reg_30__31_ ( .D(n2942), .CLK(clk), .Q(fifo_array[1291])
         );
  DFFPOSX1 fifo_array_reg_30__30_ ( .D(n2941), .CLK(clk), .Q(fifo_array[1290])
         );
  DFFPOSX1 fifo_array_reg_30__29_ ( .D(n2940), .CLK(clk), .Q(fifo_array[1289])
         );
  DFFPOSX1 fifo_array_reg_30__28_ ( .D(n2939), .CLK(clk), .Q(fifo_array[1288])
         );
  DFFPOSX1 fifo_array_reg_30__27_ ( .D(n2938), .CLK(clk), .Q(fifo_array[1287])
         );
  DFFPOSX1 fifo_array_reg_30__26_ ( .D(n2937), .CLK(clk), .Q(fifo_array[1286])
         );
  DFFPOSX1 fifo_array_reg_30__25_ ( .D(n2936), .CLK(clk), .Q(fifo_array[1285])
         );
  DFFPOSX1 fifo_array_reg_30__24_ ( .D(n2935), .CLK(clk), .Q(fifo_array[1284])
         );
  DFFPOSX1 fifo_array_reg_30__23_ ( .D(n2934), .CLK(clk), .Q(fifo_array[1283])
         );
  DFFPOSX1 fifo_array_reg_30__22_ ( .D(n2933), .CLK(clk), .Q(fifo_array[1282])
         );
  DFFPOSX1 fifo_array_reg_30__21_ ( .D(n2932), .CLK(clk), .Q(fifo_array[1281])
         );
  DFFPOSX1 fifo_array_reg_30__20_ ( .D(n2931), .CLK(clk), .Q(fifo_array[1280])
         );
  DFFPOSX1 fifo_array_reg_30__19_ ( .D(n2930), .CLK(clk), .Q(fifo_array[1279])
         );
  DFFPOSX1 fifo_array_reg_30__18_ ( .D(n2929), .CLK(clk), .Q(fifo_array[1278])
         );
  DFFPOSX1 fifo_array_reg_30__17_ ( .D(n2928), .CLK(clk), .Q(fifo_array[1277])
         );
  DFFPOSX1 fifo_array_reg_30__16_ ( .D(n2927), .CLK(clk), .Q(fifo_array[1276])
         );
  DFFPOSX1 fifo_array_reg_30__15_ ( .D(n2926), .CLK(clk), .Q(fifo_array[1275])
         );
  DFFPOSX1 fifo_array_reg_30__14_ ( .D(n2925), .CLK(clk), .Q(fifo_array[1274])
         );
  DFFPOSX1 fifo_array_reg_30__13_ ( .D(n2924), .CLK(clk), .Q(fifo_array[1273])
         );
  DFFPOSX1 fifo_array_reg_30__12_ ( .D(n2923), .CLK(clk), .Q(fifo_array[1272])
         );
  DFFPOSX1 fifo_array_reg_30__11_ ( .D(n2922), .CLK(clk), .Q(fifo_array[1271])
         );
  DFFPOSX1 fifo_array_reg_30__10_ ( .D(n2921), .CLK(clk), .Q(fifo_array[1270])
         );
  DFFPOSX1 fifo_array_reg_30__9_ ( .D(n2920), .CLK(clk), .Q(fifo_array[1269])
         );
  DFFPOSX1 fifo_array_reg_30__8_ ( .D(n2919), .CLK(clk), .Q(fifo_array[1268])
         );
  DFFPOSX1 fifo_array_reg_30__7_ ( .D(n2918), .CLK(clk), .Q(fifo_array[1267])
         );
  DFFPOSX1 fifo_array_reg_30__6_ ( .D(n2917), .CLK(clk), .Q(fifo_array[1266])
         );
  DFFPOSX1 fifo_array_reg_30__5_ ( .D(n2916), .CLK(clk), .Q(fifo_array[1265])
         );
  DFFPOSX1 fifo_array_reg_30__4_ ( .D(n2915), .CLK(clk), .Q(fifo_array[1264])
         );
  DFFPOSX1 fifo_array_reg_30__3_ ( .D(n2914), .CLK(clk), .Q(fifo_array[1263])
         );
  DFFPOSX1 fifo_array_reg_30__2_ ( .D(n2913), .CLK(clk), .Q(fifo_array[1262])
         );
  DFFPOSX1 fifo_array_reg_30__1_ ( .D(n2912), .CLK(clk), .Q(fifo_array[1261])
         );
  DFFPOSX1 fifo_array_reg_30__0_ ( .D(n2911), .CLK(clk), .Q(fifo_array[1260])
         );
  DFFPOSX1 fifo_array_reg_29__41_ ( .D(n2910), .CLK(clk), .Q(fifo_array[1259])
         );
  DFFPOSX1 fifo_array_reg_29__40_ ( .D(n2909), .CLK(clk), .Q(fifo_array[1258])
         );
  DFFPOSX1 fifo_array_reg_29__39_ ( .D(n2908), .CLK(clk), .Q(fifo_array[1257])
         );
  DFFPOSX1 fifo_array_reg_29__38_ ( .D(n2907), .CLK(clk), .Q(fifo_array[1256])
         );
  DFFPOSX1 fifo_array_reg_29__37_ ( .D(n2906), .CLK(clk), .Q(fifo_array[1255])
         );
  DFFPOSX1 fifo_array_reg_29__36_ ( .D(n2905), .CLK(clk), .Q(fifo_array[1254])
         );
  DFFPOSX1 fifo_array_reg_29__35_ ( .D(n2904), .CLK(clk), .Q(fifo_array[1253])
         );
  DFFPOSX1 fifo_array_reg_29__34_ ( .D(n2903), .CLK(clk), .Q(fifo_array[1252])
         );
  DFFPOSX1 fifo_array_reg_29__33_ ( .D(n2902), .CLK(clk), .Q(fifo_array[1251])
         );
  DFFPOSX1 fifo_array_reg_29__32_ ( .D(n2901), .CLK(clk), .Q(fifo_array[1250])
         );
  DFFPOSX1 fifo_array_reg_29__31_ ( .D(n2900), .CLK(clk), .Q(fifo_array[1249])
         );
  DFFPOSX1 fifo_array_reg_29__30_ ( .D(n2899), .CLK(clk), .Q(fifo_array[1248])
         );
  DFFPOSX1 fifo_array_reg_29__29_ ( .D(n2898), .CLK(clk), .Q(fifo_array[1247])
         );
  DFFPOSX1 fifo_array_reg_29__28_ ( .D(n2897), .CLK(clk), .Q(fifo_array[1246])
         );
  DFFPOSX1 fifo_array_reg_29__27_ ( .D(n2896), .CLK(clk), .Q(fifo_array[1245])
         );
  DFFPOSX1 fifo_array_reg_29__26_ ( .D(n2895), .CLK(clk), .Q(fifo_array[1244])
         );
  DFFPOSX1 fifo_array_reg_29__25_ ( .D(n2894), .CLK(clk), .Q(fifo_array[1243])
         );
  DFFPOSX1 fifo_array_reg_29__24_ ( .D(n2893), .CLK(clk), .Q(fifo_array[1242])
         );
  DFFPOSX1 fifo_array_reg_29__23_ ( .D(n2892), .CLK(clk), .Q(fifo_array[1241])
         );
  DFFPOSX1 fifo_array_reg_29__22_ ( .D(n2891), .CLK(clk), .Q(fifo_array[1240])
         );
  DFFPOSX1 fifo_array_reg_29__21_ ( .D(n2890), .CLK(clk), .Q(fifo_array[1239])
         );
  DFFPOSX1 fifo_array_reg_29__20_ ( .D(n2889), .CLK(clk), .Q(fifo_array[1238])
         );
  DFFPOSX1 fifo_array_reg_29__19_ ( .D(n2888), .CLK(clk), .Q(fifo_array[1237])
         );
  DFFPOSX1 fifo_array_reg_29__18_ ( .D(n2887), .CLK(clk), .Q(fifo_array[1236])
         );
  DFFPOSX1 fifo_array_reg_29__17_ ( .D(n2886), .CLK(clk), .Q(fifo_array[1235])
         );
  DFFPOSX1 fifo_array_reg_29__16_ ( .D(n2885), .CLK(clk), .Q(fifo_array[1234])
         );
  DFFPOSX1 fifo_array_reg_29__15_ ( .D(n2884), .CLK(clk), .Q(fifo_array[1233])
         );
  DFFPOSX1 fifo_array_reg_29__14_ ( .D(n2883), .CLK(clk), .Q(fifo_array[1232])
         );
  DFFPOSX1 fifo_array_reg_29__13_ ( .D(n2882), .CLK(clk), .Q(fifo_array[1231])
         );
  DFFPOSX1 fifo_array_reg_29__12_ ( .D(n2881), .CLK(clk), .Q(fifo_array[1230])
         );
  DFFPOSX1 fifo_array_reg_29__11_ ( .D(n2880), .CLK(clk), .Q(fifo_array[1229])
         );
  DFFPOSX1 fifo_array_reg_29__10_ ( .D(n2879), .CLK(clk), .Q(fifo_array[1228])
         );
  DFFPOSX1 fifo_array_reg_29__9_ ( .D(n2878), .CLK(clk), .Q(fifo_array[1227])
         );
  DFFPOSX1 fifo_array_reg_29__8_ ( .D(n2877), .CLK(clk), .Q(fifo_array[1226])
         );
  DFFPOSX1 fifo_array_reg_29__7_ ( .D(n2876), .CLK(clk), .Q(fifo_array[1225])
         );
  DFFPOSX1 fifo_array_reg_29__6_ ( .D(n2875), .CLK(clk), .Q(fifo_array[1224])
         );
  DFFPOSX1 fifo_array_reg_29__5_ ( .D(n2874), .CLK(clk), .Q(fifo_array[1223])
         );
  DFFPOSX1 fifo_array_reg_29__4_ ( .D(n2873), .CLK(clk), .Q(fifo_array[1222])
         );
  DFFPOSX1 fifo_array_reg_29__3_ ( .D(n2872), .CLK(clk), .Q(fifo_array[1221])
         );
  DFFPOSX1 fifo_array_reg_29__2_ ( .D(n2871), .CLK(clk), .Q(fifo_array[1220])
         );
  DFFPOSX1 fifo_array_reg_29__1_ ( .D(n2870), .CLK(clk), .Q(fifo_array[1219])
         );
  DFFPOSX1 fifo_array_reg_29__0_ ( .D(n2869), .CLK(clk), .Q(fifo_array[1218])
         );
  DFFPOSX1 fifo_array_reg_28__41_ ( .D(n2868), .CLK(clk), .Q(fifo_array[1217])
         );
  DFFPOSX1 fifo_array_reg_28__40_ ( .D(n2867), .CLK(clk), .Q(fifo_array[1216])
         );
  DFFPOSX1 fifo_array_reg_28__39_ ( .D(n2866), .CLK(clk), .Q(fifo_array[1215])
         );
  DFFPOSX1 fifo_array_reg_28__38_ ( .D(n2865), .CLK(clk), .Q(fifo_array[1214])
         );
  DFFPOSX1 fifo_array_reg_28__37_ ( .D(n2864), .CLK(clk), .Q(fifo_array[1213])
         );
  DFFPOSX1 fifo_array_reg_28__36_ ( .D(n2863), .CLK(clk), .Q(fifo_array[1212])
         );
  DFFPOSX1 fifo_array_reg_28__35_ ( .D(n2862), .CLK(clk), .Q(fifo_array[1211])
         );
  DFFPOSX1 fifo_array_reg_28__34_ ( .D(n2861), .CLK(clk), .Q(fifo_array[1210])
         );
  DFFPOSX1 fifo_array_reg_28__33_ ( .D(n2860), .CLK(clk), .Q(fifo_array[1209])
         );
  DFFPOSX1 fifo_array_reg_28__32_ ( .D(n2859), .CLK(clk), .Q(fifo_array[1208])
         );
  DFFPOSX1 fifo_array_reg_28__31_ ( .D(n2858), .CLK(clk), .Q(fifo_array[1207])
         );
  DFFPOSX1 fifo_array_reg_28__30_ ( .D(n2857), .CLK(clk), .Q(fifo_array[1206])
         );
  DFFPOSX1 fifo_array_reg_28__29_ ( .D(n2856), .CLK(clk), .Q(fifo_array[1205])
         );
  DFFPOSX1 fifo_array_reg_28__28_ ( .D(n2855), .CLK(clk), .Q(fifo_array[1204])
         );
  DFFPOSX1 fifo_array_reg_28__27_ ( .D(n2854), .CLK(clk), .Q(fifo_array[1203])
         );
  DFFPOSX1 fifo_array_reg_28__26_ ( .D(n2853), .CLK(clk), .Q(fifo_array[1202])
         );
  DFFPOSX1 fifo_array_reg_28__25_ ( .D(n2852), .CLK(clk), .Q(fifo_array[1201])
         );
  DFFPOSX1 fifo_array_reg_28__24_ ( .D(n2851), .CLK(clk), .Q(fifo_array[1200])
         );
  DFFPOSX1 fifo_array_reg_28__23_ ( .D(n2850), .CLK(clk), .Q(fifo_array[1199])
         );
  DFFPOSX1 fifo_array_reg_28__22_ ( .D(n2849), .CLK(clk), .Q(fifo_array[1198])
         );
  DFFPOSX1 fifo_array_reg_28__21_ ( .D(n2848), .CLK(clk), .Q(fifo_array[1197])
         );
  DFFPOSX1 fifo_array_reg_28__20_ ( .D(n2847), .CLK(clk), .Q(fifo_array[1196])
         );
  DFFPOSX1 fifo_array_reg_28__19_ ( .D(n2846), .CLK(clk), .Q(fifo_array[1195])
         );
  DFFPOSX1 fifo_array_reg_28__18_ ( .D(n2845), .CLK(clk), .Q(fifo_array[1194])
         );
  DFFPOSX1 fifo_array_reg_28__17_ ( .D(n2844), .CLK(clk), .Q(fifo_array[1193])
         );
  DFFPOSX1 fifo_array_reg_28__16_ ( .D(n2843), .CLK(clk), .Q(fifo_array[1192])
         );
  DFFPOSX1 fifo_array_reg_28__15_ ( .D(n2842), .CLK(clk), .Q(fifo_array[1191])
         );
  DFFPOSX1 fifo_array_reg_28__14_ ( .D(n2841), .CLK(clk), .Q(fifo_array[1190])
         );
  DFFPOSX1 fifo_array_reg_28__13_ ( .D(n2840), .CLK(clk), .Q(fifo_array[1189])
         );
  DFFPOSX1 fifo_array_reg_28__12_ ( .D(n2839), .CLK(clk), .Q(fifo_array[1188])
         );
  DFFPOSX1 fifo_array_reg_28__11_ ( .D(n2838), .CLK(clk), .Q(fifo_array[1187])
         );
  DFFPOSX1 fifo_array_reg_28__10_ ( .D(n2837), .CLK(clk), .Q(fifo_array[1186])
         );
  DFFPOSX1 fifo_array_reg_28__9_ ( .D(n2836), .CLK(clk), .Q(fifo_array[1185])
         );
  DFFPOSX1 fifo_array_reg_28__8_ ( .D(n2835), .CLK(clk), .Q(fifo_array[1184])
         );
  DFFPOSX1 fifo_array_reg_28__7_ ( .D(n2834), .CLK(clk), .Q(fifo_array[1183])
         );
  DFFPOSX1 fifo_array_reg_28__6_ ( .D(n2833), .CLK(clk), .Q(fifo_array[1182])
         );
  DFFPOSX1 fifo_array_reg_28__5_ ( .D(n2832), .CLK(clk), .Q(fifo_array[1181])
         );
  DFFPOSX1 fifo_array_reg_28__4_ ( .D(n2831), .CLK(clk), .Q(fifo_array[1180])
         );
  DFFPOSX1 fifo_array_reg_28__3_ ( .D(n2830), .CLK(clk), .Q(fifo_array[1179])
         );
  DFFPOSX1 fifo_array_reg_28__2_ ( .D(n2829), .CLK(clk), .Q(fifo_array[1178])
         );
  DFFPOSX1 fifo_array_reg_28__1_ ( .D(n2828), .CLK(clk), .Q(fifo_array[1177])
         );
  DFFPOSX1 fifo_array_reg_28__0_ ( .D(n2827), .CLK(clk), .Q(fifo_array[1176])
         );
  DFFPOSX1 fifo_array_reg_27__41_ ( .D(n2826), .CLK(clk), .Q(fifo_array[1175])
         );
  DFFPOSX1 fifo_array_reg_27__40_ ( .D(n2825), .CLK(clk), .Q(fifo_array[1174])
         );
  DFFPOSX1 fifo_array_reg_27__39_ ( .D(n2824), .CLK(clk), .Q(fifo_array[1173])
         );
  DFFPOSX1 fifo_array_reg_27__38_ ( .D(n2823), .CLK(clk), .Q(fifo_array[1172])
         );
  DFFPOSX1 fifo_array_reg_27__37_ ( .D(n2822), .CLK(clk), .Q(fifo_array[1171])
         );
  DFFPOSX1 fifo_array_reg_27__36_ ( .D(n2821), .CLK(clk), .Q(fifo_array[1170])
         );
  DFFPOSX1 fifo_array_reg_27__35_ ( .D(n2820), .CLK(clk), .Q(fifo_array[1169])
         );
  DFFPOSX1 fifo_array_reg_27__34_ ( .D(n2819), .CLK(clk), .Q(fifo_array[1168])
         );
  DFFPOSX1 fifo_array_reg_27__33_ ( .D(n2818), .CLK(clk), .Q(fifo_array[1167])
         );
  DFFPOSX1 fifo_array_reg_27__32_ ( .D(n2817), .CLK(clk), .Q(fifo_array[1166])
         );
  DFFPOSX1 fifo_array_reg_27__31_ ( .D(n2816), .CLK(clk), .Q(fifo_array[1165])
         );
  DFFPOSX1 fifo_array_reg_27__30_ ( .D(n2815), .CLK(clk), .Q(fifo_array[1164])
         );
  DFFPOSX1 fifo_array_reg_27__29_ ( .D(n2814), .CLK(clk), .Q(fifo_array[1163])
         );
  DFFPOSX1 fifo_array_reg_27__28_ ( .D(n2813), .CLK(clk), .Q(fifo_array[1162])
         );
  DFFPOSX1 fifo_array_reg_27__27_ ( .D(n2812), .CLK(clk), .Q(fifo_array[1161])
         );
  DFFPOSX1 fifo_array_reg_27__26_ ( .D(n2811), .CLK(clk), .Q(fifo_array[1160])
         );
  DFFPOSX1 fifo_array_reg_27__25_ ( .D(n2810), .CLK(clk), .Q(fifo_array[1159])
         );
  DFFPOSX1 fifo_array_reg_27__24_ ( .D(n2809), .CLK(clk), .Q(fifo_array[1158])
         );
  DFFPOSX1 fifo_array_reg_27__23_ ( .D(n2808), .CLK(clk), .Q(fifo_array[1157])
         );
  DFFPOSX1 fifo_array_reg_27__22_ ( .D(n2807), .CLK(clk), .Q(fifo_array[1156])
         );
  DFFPOSX1 fifo_array_reg_27__21_ ( .D(n2806), .CLK(clk), .Q(fifo_array[1155])
         );
  DFFPOSX1 fifo_array_reg_27__20_ ( .D(n2805), .CLK(clk), .Q(fifo_array[1154])
         );
  DFFPOSX1 fifo_array_reg_27__19_ ( .D(n2804), .CLK(clk), .Q(fifo_array[1153])
         );
  DFFPOSX1 fifo_array_reg_27__18_ ( .D(n2803), .CLK(clk), .Q(fifo_array[1152])
         );
  DFFPOSX1 fifo_array_reg_27__17_ ( .D(n2802), .CLK(clk), .Q(fifo_array[1151])
         );
  DFFPOSX1 fifo_array_reg_27__16_ ( .D(n2801), .CLK(clk), .Q(fifo_array[1150])
         );
  DFFPOSX1 fifo_array_reg_27__15_ ( .D(n2800), .CLK(clk), .Q(fifo_array[1149])
         );
  DFFPOSX1 fifo_array_reg_27__14_ ( .D(n2799), .CLK(clk), .Q(fifo_array[1148])
         );
  DFFPOSX1 fifo_array_reg_27__13_ ( .D(n2798), .CLK(clk), .Q(fifo_array[1147])
         );
  DFFPOSX1 fifo_array_reg_27__12_ ( .D(n2797), .CLK(clk), .Q(fifo_array[1146])
         );
  DFFPOSX1 fifo_array_reg_27__11_ ( .D(n2796), .CLK(clk), .Q(fifo_array[1145])
         );
  DFFPOSX1 fifo_array_reg_27__10_ ( .D(n2795), .CLK(clk), .Q(fifo_array[1144])
         );
  DFFPOSX1 fifo_array_reg_27__9_ ( .D(n2794), .CLK(clk), .Q(fifo_array[1143])
         );
  DFFPOSX1 fifo_array_reg_27__8_ ( .D(n2793), .CLK(clk), .Q(fifo_array[1142])
         );
  DFFPOSX1 fifo_array_reg_27__7_ ( .D(n2792), .CLK(clk), .Q(fifo_array[1141])
         );
  DFFPOSX1 fifo_array_reg_27__6_ ( .D(n2791), .CLK(clk), .Q(fifo_array[1140])
         );
  DFFPOSX1 fifo_array_reg_27__5_ ( .D(n2790), .CLK(clk), .Q(fifo_array[1139])
         );
  DFFPOSX1 fifo_array_reg_27__4_ ( .D(n2789), .CLK(clk), .Q(fifo_array[1138])
         );
  DFFPOSX1 fifo_array_reg_27__3_ ( .D(n2788), .CLK(clk), .Q(fifo_array[1137])
         );
  DFFPOSX1 fifo_array_reg_27__2_ ( .D(n2787), .CLK(clk), .Q(fifo_array[1136])
         );
  DFFPOSX1 fifo_array_reg_27__1_ ( .D(n2786), .CLK(clk), .Q(fifo_array[1135])
         );
  DFFPOSX1 fifo_array_reg_27__0_ ( .D(n2785), .CLK(clk), .Q(fifo_array[1134])
         );
  DFFPOSX1 fifo_array_reg_26__41_ ( .D(n2784), .CLK(clk), .Q(fifo_array[1133])
         );
  DFFPOSX1 fifo_array_reg_26__40_ ( .D(n2783), .CLK(clk), .Q(fifo_array[1132])
         );
  DFFPOSX1 fifo_array_reg_26__39_ ( .D(n2782), .CLK(clk), .Q(fifo_array[1131])
         );
  DFFPOSX1 fifo_array_reg_26__38_ ( .D(n2781), .CLK(clk), .Q(fifo_array[1130])
         );
  DFFPOSX1 fifo_array_reg_26__37_ ( .D(n2780), .CLK(clk), .Q(fifo_array[1129])
         );
  DFFPOSX1 fifo_array_reg_26__36_ ( .D(n2779), .CLK(clk), .Q(fifo_array[1128])
         );
  DFFPOSX1 fifo_array_reg_26__35_ ( .D(n2778), .CLK(clk), .Q(fifo_array[1127])
         );
  DFFPOSX1 fifo_array_reg_26__34_ ( .D(n2777), .CLK(clk), .Q(fifo_array[1126])
         );
  DFFPOSX1 fifo_array_reg_26__33_ ( .D(n2776), .CLK(clk), .Q(fifo_array[1125])
         );
  DFFPOSX1 fifo_array_reg_26__32_ ( .D(n2775), .CLK(clk), .Q(fifo_array[1124])
         );
  DFFPOSX1 fifo_array_reg_26__31_ ( .D(n2774), .CLK(clk), .Q(fifo_array[1123])
         );
  DFFPOSX1 fifo_array_reg_26__30_ ( .D(n2773), .CLK(clk), .Q(fifo_array[1122])
         );
  DFFPOSX1 fifo_array_reg_26__29_ ( .D(n2772), .CLK(clk), .Q(fifo_array[1121])
         );
  DFFPOSX1 fifo_array_reg_26__28_ ( .D(n2771), .CLK(clk), .Q(fifo_array[1120])
         );
  DFFPOSX1 fifo_array_reg_26__27_ ( .D(n2770), .CLK(clk), .Q(fifo_array[1119])
         );
  DFFPOSX1 fifo_array_reg_26__26_ ( .D(n2769), .CLK(clk), .Q(fifo_array[1118])
         );
  DFFPOSX1 fifo_array_reg_26__25_ ( .D(n2768), .CLK(clk), .Q(fifo_array[1117])
         );
  DFFPOSX1 fifo_array_reg_26__24_ ( .D(n2767), .CLK(clk), .Q(fifo_array[1116])
         );
  DFFPOSX1 fifo_array_reg_26__23_ ( .D(n2766), .CLK(clk), .Q(fifo_array[1115])
         );
  DFFPOSX1 fifo_array_reg_26__22_ ( .D(n2765), .CLK(clk), .Q(fifo_array[1114])
         );
  DFFPOSX1 fifo_array_reg_26__21_ ( .D(n2764), .CLK(clk), .Q(fifo_array[1113])
         );
  DFFPOSX1 fifo_array_reg_26__20_ ( .D(n2763), .CLK(clk), .Q(fifo_array[1112])
         );
  DFFPOSX1 fifo_array_reg_26__19_ ( .D(n2762), .CLK(clk), .Q(fifo_array[1111])
         );
  DFFPOSX1 fifo_array_reg_26__18_ ( .D(n2761), .CLK(clk), .Q(fifo_array[1110])
         );
  DFFPOSX1 fifo_array_reg_26__17_ ( .D(n2760), .CLK(clk), .Q(fifo_array[1109])
         );
  DFFPOSX1 fifo_array_reg_26__16_ ( .D(n2759), .CLK(clk), .Q(fifo_array[1108])
         );
  DFFPOSX1 fifo_array_reg_26__15_ ( .D(n2758), .CLK(clk), .Q(fifo_array[1107])
         );
  DFFPOSX1 fifo_array_reg_26__14_ ( .D(n2757), .CLK(clk), .Q(fifo_array[1106])
         );
  DFFPOSX1 fifo_array_reg_26__13_ ( .D(n2756), .CLK(clk), .Q(fifo_array[1105])
         );
  DFFPOSX1 fifo_array_reg_26__12_ ( .D(n2755), .CLK(clk), .Q(fifo_array[1104])
         );
  DFFPOSX1 fifo_array_reg_26__11_ ( .D(n2754), .CLK(clk), .Q(fifo_array[1103])
         );
  DFFPOSX1 fifo_array_reg_26__10_ ( .D(n2753), .CLK(clk), .Q(fifo_array[1102])
         );
  DFFPOSX1 fifo_array_reg_26__9_ ( .D(n2752), .CLK(clk), .Q(fifo_array[1101])
         );
  DFFPOSX1 fifo_array_reg_26__8_ ( .D(n2751), .CLK(clk), .Q(fifo_array[1100])
         );
  DFFPOSX1 fifo_array_reg_26__7_ ( .D(n2750), .CLK(clk), .Q(fifo_array[1099])
         );
  DFFPOSX1 fifo_array_reg_26__6_ ( .D(n2749), .CLK(clk), .Q(fifo_array[1098])
         );
  DFFPOSX1 fifo_array_reg_26__5_ ( .D(n2748), .CLK(clk), .Q(fifo_array[1097])
         );
  DFFPOSX1 fifo_array_reg_26__4_ ( .D(n2747), .CLK(clk), .Q(fifo_array[1096])
         );
  DFFPOSX1 fifo_array_reg_26__3_ ( .D(n2746), .CLK(clk), .Q(fifo_array[1095])
         );
  DFFPOSX1 fifo_array_reg_26__2_ ( .D(n2745), .CLK(clk), .Q(fifo_array[1094])
         );
  DFFPOSX1 fifo_array_reg_26__1_ ( .D(n2744), .CLK(clk), .Q(fifo_array[1093])
         );
  DFFPOSX1 fifo_array_reg_26__0_ ( .D(n2743), .CLK(clk), .Q(fifo_array[1092])
         );
  DFFPOSX1 fifo_array_reg_25__41_ ( .D(n2742), .CLK(clk), .Q(fifo_array[1091])
         );
  DFFPOSX1 fifo_array_reg_25__40_ ( .D(n2741), .CLK(clk), .Q(fifo_array[1090])
         );
  DFFPOSX1 fifo_array_reg_25__39_ ( .D(n2740), .CLK(clk), .Q(fifo_array[1089])
         );
  DFFPOSX1 fifo_array_reg_25__38_ ( .D(n2739), .CLK(clk), .Q(fifo_array[1088])
         );
  DFFPOSX1 fifo_array_reg_25__37_ ( .D(n2738), .CLK(clk), .Q(fifo_array[1087])
         );
  DFFPOSX1 fifo_array_reg_25__36_ ( .D(n2737), .CLK(clk), .Q(fifo_array[1086])
         );
  DFFPOSX1 fifo_array_reg_25__35_ ( .D(n2736), .CLK(clk), .Q(fifo_array[1085])
         );
  DFFPOSX1 fifo_array_reg_25__34_ ( .D(n2735), .CLK(clk), .Q(fifo_array[1084])
         );
  DFFPOSX1 fifo_array_reg_25__33_ ( .D(n2734), .CLK(clk), .Q(fifo_array[1083])
         );
  DFFPOSX1 fifo_array_reg_25__32_ ( .D(n2733), .CLK(clk), .Q(fifo_array[1082])
         );
  DFFPOSX1 fifo_array_reg_25__31_ ( .D(n2732), .CLK(clk), .Q(fifo_array[1081])
         );
  DFFPOSX1 fifo_array_reg_25__30_ ( .D(n2731), .CLK(clk), .Q(fifo_array[1080])
         );
  DFFPOSX1 fifo_array_reg_25__29_ ( .D(n2730), .CLK(clk), .Q(fifo_array[1079])
         );
  DFFPOSX1 fifo_array_reg_25__28_ ( .D(n2729), .CLK(clk), .Q(fifo_array[1078])
         );
  DFFPOSX1 fifo_array_reg_25__27_ ( .D(n2728), .CLK(clk), .Q(fifo_array[1077])
         );
  DFFPOSX1 fifo_array_reg_25__26_ ( .D(n2727), .CLK(clk), .Q(fifo_array[1076])
         );
  DFFPOSX1 fifo_array_reg_25__25_ ( .D(n2726), .CLK(clk), .Q(fifo_array[1075])
         );
  DFFPOSX1 fifo_array_reg_25__24_ ( .D(n2725), .CLK(clk), .Q(fifo_array[1074])
         );
  DFFPOSX1 fifo_array_reg_25__23_ ( .D(n2724), .CLK(clk), .Q(fifo_array[1073])
         );
  DFFPOSX1 fifo_array_reg_25__22_ ( .D(n2723), .CLK(clk), .Q(fifo_array[1072])
         );
  DFFPOSX1 fifo_array_reg_25__21_ ( .D(n2722), .CLK(clk), .Q(fifo_array[1071])
         );
  DFFPOSX1 fifo_array_reg_25__20_ ( .D(n2721), .CLK(clk), .Q(fifo_array[1070])
         );
  DFFPOSX1 fifo_array_reg_25__19_ ( .D(n2720), .CLK(clk), .Q(fifo_array[1069])
         );
  DFFPOSX1 fifo_array_reg_25__18_ ( .D(n2719), .CLK(clk), .Q(fifo_array[1068])
         );
  DFFPOSX1 fifo_array_reg_25__17_ ( .D(n2718), .CLK(clk), .Q(fifo_array[1067])
         );
  DFFPOSX1 fifo_array_reg_25__16_ ( .D(n2717), .CLK(clk), .Q(fifo_array[1066])
         );
  DFFPOSX1 fifo_array_reg_25__15_ ( .D(n2716), .CLK(clk), .Q(fifo_array[1065])
         );
  DFFPOSX1 fifo_array_reg_25__14_ ( .D(n2715), .CLK(clk), .Q(fifo_array[1064])
         );
  DFFPOSX1 fifo_array_reg_25__13_ ( .D(n2714), .CLK(clk), .Q(fifo_array[1063])
         );
  DFFPOSX1 fifo_array_reg_25__12_ ( .D(n2713), .CLK(clk), .Q(fifo_array[1062])
         );
  DFFPOSX1 fifo_array_reg_25__11_ ( .D(n2712), .CLK(clk), .Q(fifo_array[1061])
         );
  DFFPOSX1 fifo_array_reg_25__10_ ( .D(n2711), .CLK(clk), .Q(fifo_array[1060])
         );
  DFFPOSX1 fifo_array_reg_25__9_ ( .D(n2710), .CLK(clk), .Q(fifo_array[1059])
         );
  DFFPOSX1 fifo_array_reg_25__8_ ( .D(n2709), .CLK(clk), .Q(fifo_array[1058])
         );
  DFFPOSX1 fifo_array_reg_25__7_ ( .D(n2708), .CLK(clk), .Q(fifo_array[1057])
         );
  DFFPOSX1 fifo_array_reg_25__6_ ( .D(n2707), .CLK(clk), .Q(fifo_array[1056])
         );
  DFFPOSX1 fifo_array_reg_25__5_ ( .D(n2706), .CLK(clk), .Q(fifo_array[1055])
         );
  DFFPOSX1 fifo_array_reg_25__4_ ( .D(n2705), .CLK(clk), .Q(fifo_array[1054])
         );
  DFFPOSX1 fifo_array_reg_25__3_ ( .D(n2704), .CLK(clk), .Q(fifo_array[1053])
         );
  DFFPOSX1 fifo_array_reg_25__2_ ( .D(n2703), .CLK(clk), .Q(fifo_array[1052])
         );
  DFFPOSX1 fifo_array_reg_25__1_ ( .D(n2702), .CLK(clk), .Q(fifo_array[1051])
         );
  DFFPOSX1 fifo_array_reg_25__0_ ( .D(n2701), .CLK(clk), .Q(fifo_array[1050])
         );
  DFFPOSX1 fifo_array_reg_24__41_ ( .D(n2700), .CLK(clk), .Q(fifo_array[1049])
         );
  DFFPOSX1 fifo_array_reg_24__40_ ( .D(n2699), .CLK(clk), .Q(fifo_array[1048])
         );
  DFFPOSX1 fifo_array_reg_24__39_ ( .D(n2698), .CLK(clk), .Q(fifo_array[1047])
         );
  DFFPOSX1 fifo_array_reg_24__38_ ( .D(n2697), .CLK(clk), .Q(fifo_array[1046])
         );
  DFFPOSX1 fifo_array_reg_24__37_ ( .D(n2696), .CLK(clk), .Q(fifo_array[1045])
         );
  DFFPOSX1 fifo_array_reg_24__36_ ( .D(n2695), .CLK(clk), .Q(fifo_array[1044])
         );
  DFFPOSX1 fifo_array_reg_24__35_ ( .D(n2694), .CLK(clk), .Q(fifo_array[1043])
         );
  DFFPOSX1 fifo_array_reg_24__34_ ( .D(n2693), .CLK(clk), .Q(fifo_array[1042])
         );
  DFFPOSX1 fifo_array_reg_24__33_ ( .D(n2692), .CLK(clk), .Q(fifo_array[1041])
         );
  DFFPOSX1 fifo_array_reg_24__32_ ( .D(n2691), .CLK(clk), .Q(fifo_array[1040])
         );
  DFFPOSX1 fifo_array_reg_24__31_ ( .D(n2690), .CLK(clk), .Q(fifo_array[1039])
         );
  DFFPOSX1 fifo_array_reg_24__30_ ( .D(n2689), .CLK(clk), .Q(fifo_array[1038])
         );
  DFFPOSX1 fifo_array_reg_24__29_ ( .D(n2688), .CLK(clk), .Q(fifo_array[1037])
         );
  DFFPOSX1 fifo_array_reg_24__28_ ( .D(n2687), .CLK(clk), .Q(fifo_array[1036])
         );
  DFFPOSX1 fifo_array_reg_24__27_ ( .D(n2686), .CLK(clk), .Q(fifo_array[1035])
         );
  DFFPOSX1 fifo_array_reg_24__26_ ( .D(n2685), .CLK(clk), .Q(fifo_array[1034])
         );
  DFFPOSX1 fifo_array_reg_24__25_ ( .D(n2684), .CLK(clk), .Q(fifo_array[1033])
         );
  DFFPOSX1 fifo_array_reg_24__24_ ( .D(n2683), .CLK(clk), .Q(fifo_array[1032])
         );
  DFFPOSX1 fifo_array_reg_24__23_ ( .D(n2682), .CLK(clk), .Q(fifo_array[1031])
         );
  DFFPOSX1 fifo_array_reg_24__22_ ( .D(n2681), .CLK(clk), .Q(fifo_array[1030])
         );
  DFFPOSX1 fifo_array_reg_24__21_ ( .D(n2680), .CLK(clk), .Q(fifo_array[1029])
         );
  DFFPOSX1 fifo_array_reg_24__20_ ( .D(n2679), .CLK(clk), .Q(fifo_array[1028])
         );
  DFFPOSX1 fifo_array_reg_24__19_ ( .D(n2678), .CLK(clk), .Q(fifo_array[1027])
         );
  DFFPOSX1 fifo_array_reg_24__18_ ( .D(n2677), .CLK(clk), .Q(fifo_array[1026])
         );
  DFFPOSX1 fifo_array_reg_24__17_ ( .D(n2676), .CLK(clk), .Q(fifo_array[1025])
         );
  DFFPOSX1 fifo_array_reg_24__16_ ( .D(n2675), .CLK(clk), .Q(fifo_array[1024])
         );
  DFFPOSX1 fifo_array_reg_24__15_ ( .D(n2674), .CLK(clk), .Q(fifo_array[1023])
         );
  DFFPOSX1 fifo_array_reg_24__14_ ( .D(n2673), .CLK(clk), .Q(fifo_array[1022])
         );
  DFFPOSX1 fifo_array_reg_24__13_ ( .D(n2672), .CLK(clk), .Q(fifo_array[1021])
         );
  DFFPOSX1 fifo_array_reg_24__12_ ( .D(n2671), .CLK(clk), .Q(fifo_array[1020])
         );
  DFFPOSX1 fifo_array_reg_24__11_ ( .D(n2670), .CLK(clk), .Q(fifo_array[1019])
         );
  DFFPOSX1 fifo_array_reg_24__10_ ( .D(n2669), .CLK(clk), .Q(fifo_array[1018])
         );
  DFFPOSX1 fifo_array_reg_24__9_ ( .D(n2668), .CLK(clk), .Q(fifo_array[1017])
         );
  DFFPOSX1 fifo_array_reg_24__8_ ( .D(n2667), .CLK(clk), .Q(fifo_array[1016])
         );
  DFFPOSX1 fifo_array_reg_24__7_ ( .D(n2666), .CLK(clk), .Q(fifo_array[1015])
         );
  DFFPOSX1 fifo_array_reg_24__6_ ( .D(n2665), .CLK(clk), .Q(fifo_array[1014])
         );
  DFFPOSX1 fifo_array_reg_24__5_ ( .D(n2664), .CLK(clk), .Q(fifo_array[1013])
         );
  DFFPOSX1 fifo_array_reg_24__4_ ( .D(n2663), .CLK(clk), .Q(fifo_array[1012])
         );
  DFFPOSX1 fifo_array_reg_24__3_ ( .D(n2662), .CLK(clk), .Q(fifo_array[1011])
         );
  DFFPOSX1 fifo_array_reg_24__2_ ( .D(n2661), .CLK(clk), .Q(fifo_array[1010])
         );
  DFFPOSX1 fifo_array_reg_24__1_ ( .D(n2660), .CLK(clk), .Q(fifo_array[1009])
         );
  DFFPOSX1 fifo_array_reg_24__0_ ( .D(n2659), .CLK(clk), .Q(fifo_array[1008])
         );
  DFFPOSX1 fifo_array_reg_23__41_ ( .D(n2658), .CLK(clk), .Q(fifo_array[1007])
         );
  DFFPOSX1 fifo_array_reg_23__40_ ( .D(n2657), .CLK(clk), .Q(fifo_array[1006])
         );
  DFFPOSX1 fifo_array_reg_23__39_ ( .D(n2656), .CLK(clk), .Q(fifo_array[1005])
         );
  DFFPOSX1 fifo_array_reg_23__38_ ( .D(n2655), .CLK(clk), .Q(fifo_array[1004])
         );
  DFFPOSX1 fifo_array_reg_23__37_ ( .D(n2654), .CLK(clk), .Q(fifo_array[1003])
         );
  DFFPOSX1 fifo_array_reg_23__36_ ( .D(n2653), .CLK(clk), .Q(fifo_array[1002])
         );
  DFFPOSX1 fifo_array_reg_23__35_ ( .D(n2652), .CLK(clk), .Q(fifo_array[1001])
         );
  DFFPOSX1 fifo_array_reg_23__34_ ( .D(n2651), .CLK(clk), .Q(fifo_array[1000])
         );
  DFFPOSX1 fifo_array_reg_23__33_ ( .D(n2650), .CLK(clk), .Q(fifo_array[999])
         );
  DFFPOSX1 fifo_array_reg_23__32_ ( .D(n2649), .CLK(clk), .Q(fifo_array[998])
         );
  DFFPOSX1 fifo_array_reg_23__31_ ( .D(n2648), .CLK(clk), .Q(fifo_array[997])
         );
  DFFPOSX1 fifo_array_reg_23__30_ ( .D(n2647), .CLK(clk), .Q(fifo_array[996])
         );
  DFFPOSX1 fifo_array_reg_23__29_ ( .D(n2646), .CLK(clk), .Q(fifo_array[995])
         );
  DFFPOSX1 fifo_array_reg_23__28_ ( .D(n2645), .CLK(clk), .Q(fifo_array[994])
         );
  DFFPOSX1 fifo_array_reg_23__27_ ( .D(n2644), .CLK(clk), .Q(fifo_array[993])
         );
  DFFPOSX1 fifo_array_reg_23__26_ ( .D(n2643), .CLK(clk), .Q(fifo_array[992])
         );
  DFFPOSX1 fifo_array_reg_23__25_ ( .D(n2642), .CLK(clk), .Q(fifo_array[991])
         );
  DFFPOSX1 fifo_array_reg_23__24_ ( .D(n2641), .CLK(clk), .Q(fifo_array[990])
         );
  DFFPOSX1 fifo_array_reg_23__23_ ( .D(n2640), .CLK(clk), .Q(fifo_array[989])
         );
  DFFPOSX1 fifo_array_reg_23__22_ ( .D(n2639), .CLK(clk), .Q(fifo_array[988])
         );
  DFFPOSX1 fifo_array_reg_23__21_ ( .D(n2638), .CLK(clk), .Q(fifo_array[987])
         );
  DFFPOSX1 fifo_array_reg_23__20_ ( .D(n2637), .CLK(clk), .Q(fifo_array[986])
         );
  DFFPOSX1 fifo_array_reg_23__19_ ( .D(n2636), .CLK(clk), .Q(fifo_array[985])
         );
  DFFPOSX1 fifo_array_reg_23__18_ ( .D(n2635), .CLK(clk), .Q(fifo_array[984])
         );
  DFFPOSX1 fifo_array_reg_23__17_ ( .D(n2634), .CLK(clk), .Q(fifo_array[983])
         );
  DFFPOSX1 fifo_array_reg_23__16_ ( .D(n2633), .CLK(clk), .Q(fifo_array[982])
         );
  DFFPOSX1 fifo_array_reg_23__15_ ( .D(n2632), .CLK(clk), .Q(fifo_array[981])
         );
  DFFPOSX1 fifo_array_reg_23__14_ ( .D(n2631), .CLK(clk), .Q(fifo_array[980])
         );
  DFFPOSX1 fifo_array_reg_23__13_ ( .D(n2630), .CLK(clk), .Q(fifo_array[979])
         );
  DFFPOSX1 fifo_array_reg_23__12_ ( .D(n2629), .CLK(clk), .Q(fifo_array[978])
         );
  DFFPOSX1 fifo_array_reg_23__11_ ( .D(n2628), .CLK(clk), .Q(fifo_array[977])
         );
  DFFPOSX1 fifo_array_reg_23__10_ ( .D(n2627), .CLK(clk), .Q(fifo_array[976])
         );
  DFFPOSX1 fifo_array_reg_23__9_ ( .D(n2626), .CLK(clk), .Q(fifo_array[975])
         );
  DFFPOSX1 fifo_array_reg_23__8_ ( .D(n2625), .CLK(clk), .Q(fifo_array[974])
         );
  DFFPOSX1 fifo_array_reg_23__7_ ( .D(n2624), .CLK(clk), .Q(fifo_array[973])
         );
  DFFPOSX1 fifo_array_reg_23__6_ ( .D(n2623), .CLK(clk), .Q(fifo_array[972])
         );
  DFFPOSX1 fifo_array_reg_23__5_ ( .D(n2622), .CLK(clk), .Q(fifo_array[971])
         );
  DFFPOSX1 fifo_array_reg_23__4_ ( .D(n2621), .CLK(clk), .Q(fifo_array[970])
         );
  DFFPOSX1 fifo_array_reg_23__3_ ( .D(n2620), .CLK(clk), .Q(fifo_array[969])
         );
  DFFPOSX1 fifo_array_reg_23__2_ ( .D(n2619), .CLK(clk), .Q(fifo_array[968])
         );
  DFFPOSX1 fifo_array_reg_23__1_ ( .D(n2618), .CLK(clk), .Q(fifo_array[967])
         );
  DFFPOSX1 fifo_array_reg_23__0_ ( .D(n2617), .CLK(clk), .Q(fifo_array[966])
         );
  DFFPOSX1 fifo_array_reg_22__41_ ( .D(n2616), .CLK(clk), .Q(fifo_array[965])
         );
  DFFPOSX1 fifo_array_reg_22__40_ ( .D(n2615), .CLK(clk), .Q(fifo_array[964])
         );
  DFFPOSX1 fifo_array_reg_22__39_ ( .D(n2614), .CLK(clk), .Q(fifo_array[963])
         );
  DFFPOSX1 fifo_array_reg_22__38_ ( .D(n2613), .CLK(clk), .Q(fifo_array[962])
         );
  DFFPOSX1 fifo_array_reg_22__37_ ( .D(n2612), .CLK(clk), .Q(fifo_array[961])
         );
  DFFPOSX1 fifo_array_reg_22__36_ ( .D(n2611), .CLK(clk), .Q(fifo_array[960])
         );
  DFFPOSX1 fifo_array_reg_22__35_ ( .D(n2610), .CLK(clk), .Q(fifo_array[959])
         );
  DFFPOSX1 fifo_array_reg_22__34_ ( .D(n2609), .CLK(clk), .Q(fifo_array[958])
         );
  DFFPOSX1 fifo_array_reg_22__33_ ( .D(n2608), .CLK(clk), .Q(fifo_array[957])
         );
  DFFPOSX1 fifo_array_reg_22__32_ ( .D(n2607), .CLK(clk), .Q(fifo_array[956])
         );
  DFFPOSX1 fifo_array_reg_22__31_ ( .D(n2606), .CLK(clk), .Q(fifo_array[955])
         );
  DFFPOSX1 fifo_array_reg_22__30_ ( .D(n2605), .CLK(clk), .Q(fifo_array[954])
         );
  DFFPOSX1 fifo_array_reg_22__29_ ( .D(n2604), .CLK(clk), .Q(fifo_array[953])
         );
  DFFPOSX1 fifo_array_reg_22__28_ ( .D(n2603), .CLK(clk), .Q(fifo_array[952])
         );
  DFFPOSX1 fifo_array_reg_22__27_ ( .D(n2602), .CLK(clk), .Q(fifo_array[951])
         );
  DFFPOSX1 fifo_array_reg_22__26_ ( .D(n2601), .CLK(clk), .Q(fifo_array[950])
         );
  DFFPOSX1 fifo_array_reg_22__25_ ( .D(n2600), .CLK(clk), .Q(fifo_array[949])
         );
  DFFPOSX1 fifo_array_reg_22__24_ ( .D(n2599), .CLK(clk), .Q(fifo_array[948])
         );
  DFFPOSX1 fifo_array_reg_22__23_ ( .D(n2598), .CLK(clk), .Q(fifo_array[947])
         );
  DFFPOSX1 fifo_array_reg_22__22_ ( .D(n2597), .CLK(clk), .Q(fifo_array[946])
         );
  DFFPOSX1 fifo_array_reg_22__21_ ( .D(n2596), .CLK(clk), .Q(fifo_array[945])
         );
  DFFPOSX1 fifo_array_reg_22__20_ ( .D(n2595), .CLK(clk), .Q(fifo_array[944])
         );
  DFFPOSX1 fifo_array_reg_22__19_ ( .D(n2594), .CLK(clk), .Q(fifo_array[943])
         );
  DFFPOSX1 fifo_array_reg_22__18_ ( .D(n2593), .CLK(clk), .Q(fifo_array[942])
         );
  DFFPOSX1 fifo_array_reg_22__17_ ( .D(n2592), .CLK(clk), .Q(fifo_array[941])
         );
  DFFPOSX1 fifo_array_reg_22__16_ ( .D(n2591), .CLK(clk), .Q(fifo_array[940])
         );
  DFFPOSX1 fifo_array_reg_22__15_ ( .D(n2590), .CLK(clk), .Q(fifo_array[939])
         );
  DFFPOSX1 fifo_array_reg_22__14_ ( .D(n2589), .CLK(clk), .Q(fifo_array[938])
         );
  DFFPOSX1 fifo_array_reg_22__13_ ( .D(n2588), .CLK(clk), .Q(fifo_array[937])
         );
  DFFPOSX1 fifo_array_reg_22__12_ ( .D(n2587), .CLK(clk), .Q(fifo_array[936])
         );
  DFFPOSX1 fifo_array_reg_22__11_ ( .D(n2586), .CLK(clk), .Q(fifo_array[935])
         );
  DFFPOSX1 fifo_array_reg_22__10_ ( .D(n2585), .CLK(clk), .Q(fifo_array[934])
         );
  DFFPOSX1 fifo_array_reg_22__9_ ( .D(n2584), .CLK(clk), .Q(fifo_array[933])
         );
  DFFPOSX1 fifo_array_reg_22__8_ ( .D(n2583), .CLK(clk), .Q(fifo_array[932])
         );
  DFFPOSX1 fifo_array_reg_22__7_ ( .D(n2582), .CLK(clk), .Q(fifo_array[931])
         );
  DFFPOSX1 fifo_array_reg_22__6_ ( .D(n2581), .CLK(clk), .Q(fifo_array[930])
         );
  DFFPOSX1 fifo_array_reg_22__5_ ( .D(n2580), .CLK(clk), .Q(fifo_array[929])
         );
  DFFPOSX1 fifo_array_reg_22__4_ ( .D(n2579), .CLK(clk), .Q(fifo_array[928])
         );
  DFFPOSX1 fifo_array_reg_22__3_ ( .D(n2578), .CLK(clk), .Q(fifo_array[927])
         );
  DFFPOSX1 fifo_array_reg_22__2_ ( .D(n2577), .CLK(clk), .Q(fifo_array[926])
         );
  DFFPOSX1 fifo_array_reg_22__1_ ( .D(n2576), .CLK(clk), .Q(fifo_array[925])
         );
  DFFPOSX1 fifo_array_reg_22__0_ ( .D(n2575), .CLK(clk), .Q(fifo_array[924])
         );
  DFFPOSX1 fifo_array_reg_21__41_ ( .D(n2574), .CLK(clk), .Q(fifo_array[923])
         );
  DFFPOSX1 fifo_array_reg_21__40_ ( .D(n2573), .CLK(clk), .Q(fifo_array[922])
         );
  DFFPOSX1 fifo_array_reg_21__39_ ( .D(n2572), .CLK(clk), .Q(fifo_array[921])
         );
  DFFPOSX1 fifo_array_reg_21__38_ ( .D(n2571), .CLK(clk), .Q(fifo_array[920])
         );
  DFFPOSX1 fifo_array_reg_21__37_ ( .D(n2570), .CLK(clk), .Q(fifo_array[919])
         );
  DFFPOSX1 fifo_array_reg_21__36_ ( .D(n2569), .CLK(clk), .Q(fifo_array[918])
         );
  DFFPOSX1 fifo_array_reg_21__35_ ( .D(n2568), .CLK(clk), .Q(fifo_array[917])
         );
  DFFPOSX1 fifo_array_reg_21__34_ ( .D(n2567), .CLK(clk), .Q(fifo_array[916])
         );
  DFFPOSX1 fifo_array_reg_21__33_ ( .D(n2566), .CLK(clk), .Q(fifo_array[915])
         );
  DFFPOSX1 fifo_array_reg_21__32_ ( .D(n2565), .CLK(clk), .Q(fifo_array[914])
         );
  DFFPOSX1 fifo_array_reg_21__31_ ( .D(n2564), .CLK(clk), .Q(fifo_array[913])
         );
  DFFPOSX1 fifo_array_reg_21__30_ ( .D(n2563), .CLK(clk), .Q(fifo_array[912])
         );
  DFFPOSX1 fifo_array_reg_21__29_ ( .D(n2562), .CLK(clk), .Q(fifo_array[911])
         );
  DFFPOSX1 fifo_array_reg_21__28_ ( .D(n2561), .CLK(clk), .Q(fifo_array[910])
         );
  DFFPOSX1 fifo_array_reg_21__27_ ( .D(n2560), .CLK(clk), .Q(fifo_array[909])
         );
  DFFPOSX1 fifo_array_reg_21__26_ ( .D(n2559), .CLK(clk), .Q(fifo_array[908])
         );
  DFFPOSX1 fifo_array_reg_21__25_ ( .D(n2558), .CLK(clk), .Q(fifo_array[907])
         );
  DFFPOSX1 fifo_array_reg_21__24_ ( .D(n2557), .CLK(clk), .Q(fifo_array[906])
         );
  DFFPOSX1 fifo_array_reg_21__23_ ( .D(n2556), .CLK(clk), .Q(fifo_array[905])
         );
  DFFPOSX1 fifo_array_reg_21__22_ ( .D(n2555), .CLK(clk), .Q(fifo_array[904])
         );
  DFFPOSX1 fifo_array_reg_21__21_ ( .D(n2554), .CLK(clk), .Q(fifo_array[903])
         );
  DFFPOSX1 fifo_array_reg_21__20_ ( .D(n2553), .CLK(clk), .Q(fifo_array[902])
         );
  DFFPOSX1 fifo_array_reg_21__19_ ( .D(n2552), .CLK(clk), .Q(fifo_array[901])
         );
  DFFPOSX1 fifo_array_reg_21__18_ ( .D(n2551), .CLK(clk), .Q(fifo_array[900])
         );
  DFFPOSX1 fifo_array_reg_21__17_ ( .D(n2550), .CLK(clk), .Q(fifo_array[899])
         );
  DFFPOSX1 fifo_array_reg_21__16_ ( .D(n2549), .CLK(clk), .Q(fifo_array[898])
         );
  DFFPOSX1 fifo_array_reg_21__15_ ( .D(n2548), .CLK(clk), .Q(fifo_array[897])
         );
  DFFPOSX1 fifo_array_reg_21__14_ ( .D(n2547), .CLK(clk), .Q(fifo_array[896])
         );
  DFFPOSX1 fifo_array_reg_21__13_ ( .D(n2546), .CLK(clk), .Q(fifo_array[895])
         );
  DFFPOSX1 fifo_array_reg_21__12_ ( .D(n2545), .CLK(clk), .Q(fifo_array[894])
         );
  DFFPOSX1 fifo_array_reg_21__11_ ( .D(n2544), .CLK(clk), .Q(fifo_array[893])
         );
  DFFPOSX1 fifo_array_reg_21__10_ ( .D(n2543), .CLK(clk), .Q(fifo_array[892])
         );
  DFFPOSX1 fifo_array_reg_21__9_ ( .D(n2542), .CLK(clk), .Q(fifo_array[891])
         );
  DFFPOSX1 fifo_array_reg_21__8_ ( .D(n2541), .CLK(clk), .Q(fifo_array[890])
         );
  DFFPOSX1 fifo_array_reg_21__7_ ( .D(n2540), .CLK(clk), .Q(fifo_array[889])
         );
  DFFPOSX1 fifo_array_reg_21__6_ ( .D(n2539), .CLK(clk), .Q(fifo_array[888])
         );
  DFFPOSX1 fifo_array_reg_21__5_ ( .D(n2538), .CLK(clk), .Q(fifo_array[887])
         );
  DFFPOSX1 fifo_array_reg_21__4_ ( .D(n2537), .CLK(clk), .Q(fifo_array[886])
         );
  DFFPOSX1 fifo_array_reg_21__3_ ( .D(n2536), .CLK(clk), .Q(fifo_array[885])
         );
  DFFPOSX1 fifo_array_reg_21__2_ ( .D(n2535), .CLK(clk), .Q(fifo_array[884])
         );
  DFFPOSX1 fifo_array_reg_21__1_ ( .D(n2534), .CLK(clk), .Q(fifo_array[883])
         );
  DFFPOSX1 fifo_array_reg_21__0_ ( .D(n2533), .CLK(clk), .Q(fifo_array[882])
         );
  DFFPOSX1 fifo_array_reg_20__41_ ( .D(n2532), .CLK(clk), .Q(fifo_array[881])
         );
  DFFPOSX1 fifo_array_reg_20__40_ ( .D(n2531), .CLK(clk), .Q(fifo_array[880])
         );
  DFFPOSX1 fifo_array_reg_20__39_ ( .D(n2530), .CLK(clk), .Q(fifo_array[879])
         );
  DFFPOSX1 fifo_array_reg_20__38_ ( .D(n2529), .CLK(clk), .Q(fifo_array[878])
         );
  DFFPOSX1 fifo_array_reg_20__37_ ( .D(n2528), .CLK(clk), .Q(fifo_array[877])
         );
  DFFPOSX1 fifo_array_reg_20__36_ ( .D(n2527), .CLK(clk), .Q(fifo_array[876])
         );
  DFFPOSX1 fifo_array_reg_20__35_ ( .D(n2526), .CLK(clk), .Q(fifo_array[875])
         );
  DFFPOSX1 fifo_array_reg_20__34_ ( .D(n2525), .CLK(clk), .Q(fifo_array[874])
         );
  DFFPOSX1 fifo_array_reg_20__33_ ( .D(n2524), .CLK(clk), .Q(fifo_array[873])
         );
  DFFPOSX1 fifo_array_reg_20__32_ ( .D(n2523), .CLK(clk), .Q(fifo_array[872])
         );
  DFFPOSX1 fifo_array_reg_20__31_ ( .D(n2522), .CLK(clk), .Q(fifo_array[871])
         );
  DFFPOSX1 fifo_array_reg_20__30_ ( .D(n2521), .CLK(clk), .Q(fifo_array[870])
         );
  DFFPOSX1 fifo_array_reg_20__29_ ( .D(n2520), .CLK(clk), .Q(fifo_array[869])
         );
  DFFPOSX1 fifo_array_reg_20__28_ ( .D(n2519), .CLK(clk), .Q(fifo_array[868])
         );
  DFFPOSX1 fifo_array_reg_20__27_ ( .D(n2518), .CLK(clk), .Q(fifo_array[867])
         );
  DFFPOSX1 fifo_array_reg_20__26_ ( .D(n2517), .CLK(clk), .Q(fifo_array[866])
         );
  DFFPOSX1 fifo_array_reg_20__25_ ( .D(n2516), .CLK(clk), .Q(fifo_array[865])
         );
  DFFPOSX1 fifo_array_reg_20__24_ ( .D(n2515), .CLK(clk), .Q(fifo_array[864])
         );
  DFFPOSX1 fifo_array_reg_20__23_ ( .D(n2514), .CLK(clk), .Q(fifo_array[863])
         );
  DFFPOSX1 fifo_array_reg_20__22_ ( .D(n2513), .CLK(clk), .Q(fifo_array[862])
         );
  DFFPOSX1 fifo_array_reg_20__21_ ( .D(n2512), .CLK(clk), .Q(fifo_array[861])
         );
  DFFPOSX1 fifo_array_reg_20__20_ ( .D(n2511), .CLK(clk), .Q(fifo_array[860])
         );
  DFFPOSX1 fifo_array_reg_20__19_ ( .D(n2510), .CLK(clk), .Q(fifo_array[859])
         );
  DFFPOSX1 fifo_array_reg_20__18_ ( .D(n2509), .CLK(clk), .Q(fifo_array[858])
         );
  DFFPOSX1 fifo_array_reg_20__17_ ( .D(n2508), .CLK(clk), .Q(fifo_array[857])
         );
  DFFPOSX1 fifo_array_reg_20__16_ ( .D(n2507), .CLK(clk), .Q(fifo_array[856])
         );
  DFFPOSX1 fifo_array_reg_20__15_ ( .D(n2506), .CLK(clk), .Q(fifo_array[855])
         );
  DFFPOSX1 fifo_array_reg_20__14_ ( .D(n2505), .CLK(clk), .Q(fifo_array[854])
         );
  DFFPOSX1 fifo_array_reg_20__13_ ( .D(n2504), .CLK(clk), .Q(fifo_array[853])
         );
  DFFPOSX1 fifo_array_reg_20__12_ ( .D(n2503), .CLK(clk), .Q(fifo_array[852])
         );
  DFFPOSX1 fifo_array_reg_20__11_ ( .D(n2502), .CLK(clk), .Q(fifo_array[851])
         );
  DFFPOSX1 fifo_array_reg_20__10_ ( .D(n2501), .CLK(clk), .Q(fifo_array[850])
         );
  DFFPOSX1 fifo_array_reg_20__9_ ( .D(n2500), .CLK(clk), .Q(fifo_array[849])
         );
  DFFPOSX1 fifo_array_reg_20__8_ ( .D(n2499), .CLK(clk), .Q(fifo_array[848])
         );
  DFFPOSX1 fifo_array_reg_20__7_ ( .D(n2498), .CLK(clk), .Q(fifo_array[847])
         );
  DFFPOSX1 fifo_array_reg_20__6_ ( .D(n2497), .CLK(clk), .Q(fifo_array[846])
         );
  DFFPOSX1 fifo_array_reg_20__5_ ( .D(n2496), .CLK(clk), .Q(fifo_array[845])
         );
  DFFPOSX1 fifo_array_reg_20__4_ ( .D(n2495), .CLK(clk), .Q(fifo_array[844])
         );
  DFFPOSX1 fifo_array_reg_20__3_ ( .D(n2494), .CLK(clk), .Q(fifo_array[843])
         );
  DFFPOSX1 fifo_array_reg_20__2_ ( .D(n2493), .CLK(clk), .Q(fifo_array[842])
         );
  DFFPOSX1 fifo_array_reg_20__1_ ( .D(n2492), .CLK(clk), .Q(fifo_array[841])
         );
  DFFPOSX1 fifo_array_reg_20__0_ ( .D(n2491), .CLK(clk), .Q(fifo_array[840])
         );
  DFFPOSX1 fifo_array_reg_19__41_ ( .D(n2490), .CLK(clk), .Q(fifo_array[839])
         );
  DFFPOSX1 fifo_array_reg_19__40_ ( .D(n2489), .CLK(clk), .Q(fifo_array[838])
         );
  DFFPOSX1 fifo_array_reg_19__39_ ( .D(n2488), .CLK(clk), .Q(fifo_array[837])
         );
  DFFPOSX1 fifo_array_reg_19__38_ ( .D(n2487), .CLK(clk), .Q(fifo_array[836])
         );
  DFFPOSX1 fifo_array_reg_19__37_ ( .D(n2486), .CLK(clk), .Q(fifo_array[835])
         );
  DFFPOSX1 fifo_array_reg_19__36_ ( .D(n2485), .CLK(clk), .Q(fifo_array[834])
         );
  DFFPOSX1 fifo_array_reg_19__35_ ( .D(n2484), .CLK(clk), .Q(fifo_array[833])
         );
  DFFPOSX1 fifo_array_reg_19__34_ ( .D(n2483), .CLK(clk), .Q(fifo_array[832])
         );
  DFFPOSX1 fifo_array_reg_19__33_ ( .D(n2482), .CLK(clk), .Q(fifo_array[831])
         );
  DFFPOSX1 fifo_array_reg_19__32_ ( .D(n2481), .CLK(clk), .Q(fifo_array[830])
         );
  DFFPOSX1 fifo_array_reg_19__31_ ( .D(n2480), .CLK(clk), .Q(fifo_array[829])
         );
  DFFPOSX1 fifo_array_reg_19__30_ ( .D(n2479), .CLK(clk), .Q(fifo_array[828])
         );
  DFFPOSX1 fifo_array_reg_19__29_ ( .D(n2478), .CLK(clk), .Q(fifo_array[827])
         );
  DFFPOSX1 fifo_array_reg_19__28_ ( .D(n2477), .CLK(clk), .Q(fifo_array[826])
         );
  DFFPOSX1 fifo_array_reg_19__27_ ( .D(n2476), .CLK(clk), .Q(fifo_array[825])
         );
  DFFPOSX1 fifo_array_reg_19__26_ ( .D(n2475), .CLK(clk), .Q(fifo_array[824])
         );
  DFFPOSX1 fifo_array_reg_19__25_ ( .D(n2474), .CLK(clk), .Q(fifo_array[823])
         );
  DFFPOSX1 fifo_array_reg_19__24_ ( .D(n2473), .CLK(clk), .Q(fifo_array[822])
         );
  DFFPOSX1 fifo_array_reg_19__23_ ( .D(n2472), .CLK(clk), .Q(fifo_array[821])
         );
  DFFPOSX1 fifo_array_reg_19__22_ ( .D(n2471), .CLK(clk), .Q(fifo_array[820])
         );
  DFFPOSX1 fifo_array_reg_19__21_ ( .D(n2470), .CLK(clk), .Q(fifo_array[819])
         );
  DFFPOSX1 fifo_array_reg_19__20_ ( .D(n2469), .CLK(clk), .Q(fifo_array[818])
         );
  DFFPOSX1 fifo_array_reg_19__19_ ( .D(n2468), .CLK(clk), .Q(fifo_array[817])
         );
  DFFPOSX1 fifo_array_reg_19__18_ ( .D(n2467), .CLK(clk), .Q(fifo_array[816])
         );
  DFFPOSX1 fifo_array_reg_19__17_ ( .D(n2466), .CLK(clk), .Q(fifo_array[815])
         );
  DFFPOSX1 fifo_array_reg_19__16_ ( .D(n2465), .CLK(clk), .Q(fifo_array[814])
         );
  DFFPOSX1 fifo_array_reg_19__15_ ( .D(n2464), .CLK(clk), .Q(fifo_array[813])
         );
  DFFPOSX1 fifo_array_reg_19__14_ ( .D(n2463), .CLK(clk), .Q(fifo_array[812])
         );
  DFFPOSX1 fifo_array_reg_19__13_ ( .D(n2462), .CLK(clk), .Q(fifo_array[811])
         );
  DFFPOSX1 fifo_array_reg_19__12_ ( .D(n2461), .CLK(clk), .Q(fifo_array[810])
         );
  DFFPOSX1 fifo_array_reg_19__11_ ( .D(n2460), .CLK(clk), .Q(fifo_array[809])
         );
  DFFPOSX1 fifo_array_reg_19__10_ ( .D(n2459), .CLK(clk), .Q(fifo_array[808])
         );
  DFFPOSX1 fifo_array_reg_19__9_ ( .D(n2458), .CLK(clk), .Q(fifo_array[807])
         );
  DFFPOSX1 fifo_array_reg_19__8_ ( .D(n2457), .CLK(clk), .Q(fifo_array[806])
         );
  DFFPOSX1 fifo_array_reg_19__7_ ( .D(n2456), .CLK(clk), .Q(fifo_array[805])
         );
  DFFPOSX1 fifo_array_reg_19__6_ ( .D(n2455), .CLK(clk), .Q(fifo_array[804])
         );
  DFFPOSX1 fifo_array_reg_19__5_ ( .D(n2454), .CLK(clk), .Q(fifo_array[803])
         );
  DFFPOSX1 fifo_array_reg_19__4_ ( .D(n2453), .CLK(clk), .Q(fifo_array[802])
         );
  DFFPOSX1 fifo_array_reg_19__3_ ( .D(n2452), .CLK(clk), .Q(fifo_array[801])
         );
  DFFPOSX1 fifo_array_reg_19__2_ ( .D(n2451), .CLK(clk), .Q(fifo_array[800])
         );
  DFFPOSX1 fifo_array_reg_19__1_ ( .D(n2450), .CLK(clk), .Q(fifo_array[799])
         );
  DFFPOSX1 fifo_array_reg_19__0_ ( .D(n2449), .CLK(clk), .Q(fifo_array[798])
         );
  DFFPOSX1 fifo_array_reg_18__41_ ( .D(n2448), .CLK(clk), .Q(fifo_array[797])
         );
  DFFPOSX1 fifo_array_reg_18__40_ ( .D(n2447), .CLK(clk), .Q(fifo_array[796])
         );
  DFFPOSX1 fifo_array_reg_18__39_ ( .D(n2446), .CLK(clk), .Q(fifo_array[795])
         );
  DFFPOSX1 fifo_array_reg_18__38_ ( .D(n2445), .CLK(clk), .Q(fifo_array[794])
         );
  DFFPOSX1 fifo_array_reg_18__37_ ( .D(n2444), .CLK(clk), .Q(fifo_array[793])
         );
  DFFPOSX1 fifo_array_reg_18__36_ ( .D(n2443), .CLK(clk), .Q(fifo_array[792])
         );
  DFFPOSX1 fifo_array_reg_18__35_ ( .D(n2442), .CLK(clk), .Q(fifo_array[791])
         );
  DFFPOSX1 fifo_array_reg_18__34_ ( .D(n2441), .CLK(clk), .Q(fifo_array[790])
         );
  DFFPOSX1 fifo_array_reg_18__33_ ( .D(n2440), .CLK(clk), .Q(fifo_array[789])
         );
  DFFPOSX1 fifo_array_reg_18__32_ ( .D(n2439), .CLK(clk), .Q(fifo_array[788])
         );
  DFFPOSX1 fifo_array_reg_18__31_ ( .D(n2438), .CLK(clk), .Q(fifo_array[787])
         );
  DFFPOSX1 fifo_array_reg_18__30_ ( .D(n2437), .CLK(clk), .Q(fifo_array[786])
         );
  DFFPOSX1 fifo_array_reg_18__29_ ( .D(n2436), .CLK(clk), .Q(fifo_array[785])
         );
  DFFPOSX1 fifo_array_reg_18__28_ ( .D(n2435), .CLK(clk), .Q(fifo_array[784])
         );
  DFFPOSX1 fifo_array_reg_18__27_ ( .D(n2434), .CLK(clk), .Q(fifo_array[783])
         );
  DFFPOSX1 fifo_array_reg_18__26_ ( .D(n2433), .CLK(clk), .Q(fifo_array[782])
         );
  DFFPOSX1 fifo_array_reg_18__25_ ( .D(n2432), .CLK(clk), .Q(fifo_array[781])
         );
  DFFPOSX1 fifo_array_reg_18__24_ ( .D(n2431), .CLK(clk), .Q(fifo_array[780])
         );
  DFFPOSX1 fifo_array_reg_18__23_ ( .D(n2430), .CLK(clk), .Q(fifo_array[779])
         );
  DFFPOSX1 fifo_array_reg_18__22_ ( .D(n2429), .CLK(clk), .Q(fifo_array[778])
         );
  DFFPOSX1 fifo_array_reg_18__21_ ( .D(n2428), .CLK(clk), .Q(fifo_array[777])
         );
  DFFPOSX1 fifo_array_reg_18__20_ ( .D(n2427), .CLK(clk), .Q(fifo_array[776])
         );
  DFFPOSX1 fifo_array_reg_18__19_ ( .D(n2426), .CLK(clk), .Q(fifo_array[775])
         );
  DFFPOSX1 fifo_array_reg_18__18_ ( .D(n2425), .CLK(clk), .Q(fifo_array[774])
         );
  DFFPOSX1 fifo_array_reg_18__17_ ( .D(n2424), .CLK(clk), .Q(fifo_array[773])
         );
  DFFPOSX1 fifo_array_reg_18__16_ ( .D(n2423), .CLK(clk), .Q(fifo_array[772])
         );
  DFFPOSX1 fifo_array_reg_18__15_ ( .D(n2422), .CLK(clk), .Q(fifo_array[771])
         );
  DFFPOSX1 fifo_array_reg_18__14_ ( .D(n2421), .CLK(clk), .Q(fifo_array[770])
         );
  DFFPOSX1 fifo_array_reg_18__13_ ( .D(n2420), .CLK(clk), .Q(fifo_array[769])
         );
  DFFPOSX1 fifo_array_reg_18__12_ ( .D(n2419), .CLK(clk), .Q(fifo_array[768])
         );
  DFFPOSX1 fifo_array_reg_18__11_ ( .D(n2418), .CLK(clk), .Q(fifo_array[767])
         );
  DFFPOSX1 fifo_array_reg_18__10_ ( .D(n2417), .CLK(clk), .Q(fifo_array[766])
         );
  DFFPOSX1 fifo_array_reg_18__9_ ( .D(n2416), .CLK(clk), .Q(fifo_array[765])
         );
  DFFPOSX1 fifo_array_reg_18__8_ ( .D(n2415), .CLK(clk), .Q(fifo_array[764])
         );
  DFFPOSX1 fifo_array_reg_18__7_ ( .D(n2414), .CLK(clk), .Q(fifo_array[763])
         );
  DFFPOSX1 fifo_array_reg_18__6_ ( .D(n2413), .CLK(clk), .Q(fifo_array[762])
         );
  DFFPOSX1 fifo_array_reg_18__5_ ( .D(n2412), .CLK(clk), .Q(fifo_array[761])
         );
  DFFPOSX1 fifo_array_reg_18__4_ ( .D(n2411), .CLK(clk), .Q(fifo_array[760])
         );
  DFFPOSX1 fifo_array_reg_18__3_ ( .D(n2410), .CLK(clk), .Q(fifo_array[759])
         );
  DFFPOSX1 fifo_array_reg_18__2_ ( .D(n2409), .CLK(clk), .Q(fifo_array[758])
         );
  DFFPOSX1 fifo_array_reg_18__1_ ( .D(n2408), .CLK(clk), .Q(fifo_array[757])
         );
  DFFPOSX1 fifo_array_reg_18__0_ ( .D(n2407), .CLK(clk), .Q(fifo_array[756])
         );
  DFFPOSX1 fifo_array_reg_17__41_ ( .D(n2406), .CLK(clk), .Q(fifo_array[755])
         );
  DFFPOSX1 fifo_array_reg_17__40_ ( .D(n2405), .CLK(clk), .Q(fifo_array[754])
         );
  DFFPOSX1 fifo_array_reg_17__39_ ( .D(n2404), .CLK(clk), .Q(fifo_array[753])
         );
  DFFPOSX1 fifo_array_reg_17__38_ ( .D(n2403), .CLK(clk), .Q(fifo_array[752])
         );
  DFFPOSX1 fifo_array_reg_17__37_ ( .D(n2402), .CLK(clk), .Q(fifo_array[751])
         );
  DFFPOSX1 fifo_array_reg_17__36_ ( .D(n2401), .CLK(clk), .Q(fifo_array[750])
         );
  DFFPOSX1 fifo_array_reg_17__35_ ( .D(n2400), .CLK(clk), .Q(fifo_array[749])
         );
  DFFPOSX1 fifo_array_reg_17__34_ ( .D(n2399), .CLK(clk), .Q(fifo_array[748])
         );
  DFFPOSX1 fifo_array_reg_17__33_ ( .D(n2398), .CLK(clk), .Q(fifo_array[747])
         );
  DFFPOSX1 fifo_array_reg_17__32_ ( .D(n2397), .CLK(clk), .Q(fifo_array[746])
         );
  DFFPOSX1 fifo_array_reg_17__31_ ( .D(n2396), .CLK(clk), .Q(fifo_array[745])
         );
  DFFPOSX1 fifo_array_reg_17__30_ ( .D(n2395), .CLK(clk), .Q(fifo_array[744])
         );
  DFFPOSX1 fifo_array_reg_17__29_ ( .D(n2394), .CLK(clk), .Q(fifo_array[743])
         );
  DFFPOSX1 fifo_array_reg_17__28_ ( .D(n2393), .CLK(clk), .Q(fifo_array[742])
         );
  DFFPOSX1 fifo_array_reg_17__27_ ( .D(n2392), .CLK(clk), .Q(fifo_array[741])
         );
  DFFPOSX1 fifo_array_reg_17__26_ ( .D(n2391), .CLK(clk), .Q(fifo_array[740])
         );
  DFFPOSX1 fifo_array_reg_17__25_ ( .D(n2390), .CLK(clk), .Q(fifo_array[739])
         );
  DFFPOSX1 fifo_array_reg_17__24_ ( .D(n2389), .CLK(clk), .Q(fifo_array[738])
         );
  DFFPOSX1 fifo_array_reg_17__23_ ( .D(n2388), .CLK(clk), .Q(fifo_array[737])
         );
  DFFPOSX1 fifo_array_reg_17__22_ ( .D(n2387), .CLK(clk), .Q(fifo_array[736])
         );
  DFFPOSX1 fifo_array_reg_17__21_ ( .D(n2386), .CLK(clk), .Q(fifo_array[735])
         );
  DFFPOSX1 fifo_array_reg_17__20_ ( .D(n2385), .CLK(clk), .Q(fifo_array[734])
         );
  DFFPOSX1 fifo_array_reg_17__19_ ( .D(n2384), .CLK(clk), .Q(fifo_array[733])
         );
  DFFPOSX1 fifo_array_reg_17__18_ ( .D(n2383), .CLK(clk), .Q(fifo_array[732])
         );
  DFFPOSX1 fifo_array_reg_17__17_ ( .D(n2382), .CLK(clk), .Q(fifo_array[731])
         );
  DFFPOSX1 fifo_array_reg_17__16_ ( .D(n2381), .CLK(clk), .Q(fifo_array[730])
         );
  DFFPOSX1 fifo_array_reg_17__15_ ( .D(n2380), .CLK(clk), .Q(fifo_array[729])
         );
  DFFPOSX1 fifo_array_reg_17__14_ ( .D(n2379), .CLK(clk), .Q(fifo_array[728])
         );
  DFFPOSX1 fifo_array_reg_17__13_ ( .D(n2378), .CLK(clk), .Q(fifo_array[727])
         );
  DFFPOSX1 fifo_array_reg_17__12_ ( .D(n2377), .CLK(clk), .Q(fifo_array[726])
         );
  DFFPOSX1 fifo_array_reg_17__11_ ( .D(n2376), .CLK(clk), .Q(fifo_array[725])
         );
  DFFPOSX1 fifo_array_reg_17__10_ ( .D(n2375), .CLK(clk), .Q(fifo_array[724])
         );
  DFFPOSX1 fifo_array_reg_17__9_ ( .D(n2374), .CLK(clk), .Q(fifo_array[723])
         );
  DFFPOSX1 fifo_array_reg_17__8_ ( .D(n2373), .CLK(clk), .Q(fifo_array[722])
         );
  DFFPOSX1 fifo_array_reg_17__7_ ( .D(n2372), .CLK(clk), .Q(fifo_array[721])
         );
  DFFPOSX1 fifo_array_reg_17__6_ ( .D(n2371), .CLK(clk), .Q(fifo_array[720])
         );
  DFFPOSX1 fifo_array_reg_17__5_ ( .D(n2370), .CLK(clk), .Q(fifo_array[719])
         );
  DFFPOSX1 fifo_array_reg_17__4_ ( .D(n2369), .CLK(clk), .Q(fifo_array[718])
         );
  DFFPOSX1 fifo_array_reg_17__3_ ( .D(n2368), .CLK(clk), .Q(fifo_array[717])
         );
  DFFPOSX1 fifo_array_reg_17__2_ ( .D(n2367), .CLK(clk), .Q(fifo_array[716])
         );
  DFFPOSX1 fifo_array_reg_17__1_ ( .D(n2366), .CLK(clk), .Q(fifo_array[715])
         );
  DFFPOSX1 fifo_array_reg_17__0_ ( .D(n2365), .CLK(clk), .Q(fifo_array[714])
         );
  DFFPOSX1 fifo_array_reg_16__41_ ( .D(n2364), .CLK(clk), .Q(fifo_array[713])
         );
  DFFPOSX1 fifo_array_reg_16__40_ ( .D(n2363), .CLK(clk), .Q(fifo_array[712])
         );
  DFFPOSX1 fifo_array_reg_16__39_ ( .D(n2362), .CLK(clk), .Q(fifo_array[711])
         );
  DFFPOSX1 fifo_array_reg_16__38_ ( .D(n2361), .CLK(clk), .Q(fifo_array[710])
         );
  DFFPOSX1 fifo_array_reg_16__37_ ( .D(n2360), .CLK(clk), .Q(fifo_array[709])
         );
  DFFPOSX1 fifo_array_reg_16__36_ ( .D(n2359), .CLK(clk), .Q(fifo_array[708])
         );
  DFFPOSX1 fifo_array_reg_16__35_ ( .D(n2358), .CLK(clk), .Q(fifo_array[707])
         );
  DFFPOSX1 fifo_array_reg_16__34_ ( .D(n2357), .CLK(clk), .Q(fifo_array[706])
         );
  DFFPOSX1 fifo_array_reg_16__33_ ( .D(n2356), .CLK(clk), .Q(fifo_array[705])
         );
  DFFPOSX1 fifo_array_reg_16__32_ ( .D(n2355), .CLK(clk), .Q(fifo_array[704])
         );
  DFFPOSX1 fifo_array_reg_16__31_ ( .D(n2354), .CLK(clk), .Q(fifo_array[703])
         );
  DFFPOSX1 fifo_array_reg_16__30_ ( .D(n2353), .CLK(clk), .Q(fifo_array[702])
         );
  DFFPOSX1 fifo_array_reg_16__29_ ( .D(n2352), .CLK(clk), .Q(fifo_array[701])
         );
  DFFPOSX1 fifo_array_reg_16__28_ ( .D(n2351), .CLK(clk), .Q(fifo_array[700])
         );
  DFFPOSX1 fifo_array_reg_16__27_ ( .D(n2350), .CLK(clk), .Q(fifo_array[699])
         );
  DFFPOSX1 fifo_array_reg_16__26_ ( .D(n2349), .CLK(clk), .Q(fifo_array[698])
         );
  DFFPOSX1 fifo_array_reg_16__25_ ( .D(n2348), .CLK(clk), .Q(fifo_array[697])
         );
  DFFPOSX1 fifo_array_reg_16__24_ ( .D(n2347), .CLK(clk), .Q(fifo_array[696])
         );
  DFFPOSX1 fifo_array_reg_16__23_ ( .D(n2346), .CLK(clk), .Q(fifo_array[695])
         );
  DFFPOSX1 fifo_array_reg_16__22_ ( .D(n2345), .CLK(clk), .Q(fifo_array[694])
         );
  DFFPOSX1 fifo_array_reg_16__21_ ( .D(n2344), .CLK(clk), .Q(fifo_array[693])
         );
  DFFPOSX1 fifo_array_reg_16__20_ ( .D(n2343), .CLK(clk), .Q(fifo_array[692])
         );
  DFFPOSX1 fifo_array_reg_16__19_ ( .D(n2342), .CLK(clk), .Q(fifo_array[691])
         );
  DFFPOSX1 fifo_array_reg_16__18_ ( .D(n2341), .CLK(clk), .Q(fifo_array[690])
         );
  DFFPOSX1 fifo_array_reg_16__17_ ( .D(n2340), .CLK(clk), .Q(fifo_array[689])
         );
  DFFPOSX1 fifo_array_reg_16__16_ ( .D(n2339), .CLK(clk), .Q(fifo_array[688])
         );
  DFFPOSX1 fifo_array_reg_16__15_ ( .D(n2338), .CLK(clk), .Q(fifo_array[687])
         );
  DFFPOSX1 fifo_array_reg_16__14_ ( .D(n2337), .CLK(clk), .Q(fifo_array[686])
         );
  DFFPOSX1 fifo_array_reg_16__13_ ( .D(n2336), .CLK(clk), .Q(fifo_array[685])
         );
  DFFPOSX1 fifo_array_reg_16__12_ ( .D(n2335), .CLK(clk), .Q(fifo_array[684])
         );
  DFFPOSX1 fifo_array_reg_16__11_ ( .D(n2334), .CLK(clk), .Q(fifo_array[683])
         );
  DFFPOSX1 fifo_array_reg_16__10_ ( .D(n2333), .CLK(clk), .Q(fifo_array[682])
         );
  DFFPOSX1 fifo_array_reg_16__9_ ( .D(n2332), .CLK(clk), .Q(fifo_array[681])
         );
  DFFPOSX1 fifo_array_reg_16__8_ ( .D(n2331), .CLK(clk), .Q(fifo_array[680])
         );
  DFFPOSX1 fifo_array_reg_16__7_ ( .D(n2330), .CLK(clk), .Q(fifo_array[679])
         );
  DFFPOSX1 fifo_array_reg_16__6_ ( .D(n2329), .CLK(clk), .Q(fifo_array[678])
         );
  DFFPOSX1 fifo_array_reg_16__5_ ( .D(n2328), .CLK(clk), .Q(fifo_array[677])
         );
  DFFPOSX1 fifo_array_reg_16__4_ ( .D(n2327), .CLK(clk), .Q(fifo_array[676])
         );
  DFFPOSX1 fifo_array_reg_16__3_ ( .D(n2326), .CLK(clk), .Q(fifo_array[675])
         );
  DFFPOSX1 fifo_array_reg_16__2_ ( .D(n2325), .CLK(clk), .Q(fifo_array[674])
         );
  DFFPOSX1 fifo_array_reg_16__1_ ( .D(n2324), .CLK(clk), .Q(fifo_array[673])
         );
  DFFPOSX1 fifo_array_reg_16__0_ ( .D(n2323), .CLK(clk), .Q(fifo_array[672])
         );
  DFFPOSX1 fifo_array_reg_15__41_ ( .D(n2322), .CLK(clk), .Q(fifo_array[671])
         );
  DFFPOSX1 fifo_array_reg_15__40_ ( .D(n2321), .CLK(clk), .Q(fifo_array[670])
         );
  DFFPOSX1 fifo_array_reg_15__39_ ( .D(n2320), .CLK(clk), .Q(fifo_array[669])
         );
  DFFPOSX1 fifo_array_reg_15__38_ ( .D(n2319), .CLK(clk), .Q(fifo_array[668])
         );
  DFFPOSX1 fifo_array_reg_15__37_ ( .D(n2318), .CLK(clk), .Q(fifo_array[667])
         );
  DFFPOSX1 fifo_array_reg_15__36_ ( .D(n2317), .CLK(clk), .Q(fifo_array[666])
         );
  DFFPOSX1 fifo_array_reg_15__35_ ( .D(n2316), .CLK(clk), .Q(fifo_array[665])
         );
  DFFPOSX1 fifo_array_reg_15__34_ ( .D(n2315), .CLK(clk), .Q(fifo_array[664])
         );
  DFFPOSX1 fifo_array_reg_15__33_ ( .D(n2314), .CLK(clk), .Q(fifo_array[663])
         );
  DFFPOSX1 fifo_array_reg_15__32_ ( .D(n2313), .CLK(clk), .Q(fifo_array[662])
         );
  DFFPOSX1 fifo_array_reg_15__31_ ( .D(n2312), .CLK(clk), .Q(fifo_array[661])
         );
  DFFPOSX1 fifo_array_reg_15__30_ ( .D(n2311), .CLK(clk), .Q(fifo_array[660])
         );
  DFFPOSX1 fifo_array_reg_15__29_ ( .D(n2310), .CLK(clk), .Q(fifo_array[659])
         );
  DFFPOSX1 fifo_array_reg_15__28_ ( .D(n2309), .CLK(clk), .Q(fifo_array[658])
         );
  DFFPOSX1 fifo_array_reg_15__27_ ( .D(n2308), .CLK(clk), .Q(fifo_array[657])
         );
  DFFPOSX1 fifo_array_reg_15__26_ ( .D(n2307), .CLK(clk), .Q(fifo_array[656])
         );
  DFFPOSX1 fifo_array_reg_15__25_ ( .D(n2306), .CLK(clk), .Q(fifo_array[655])
         );
  DFFPOSX1 fifo_array_reg_15__24_ ( .D(n2305), .CLK(clk), .Q(fifo_array[654])
         );
  DFFPOSX1 fifo_array_reg_15__23_ ( .D(n2304), .CLK(clk), .Q(fifo_array[653])
         );
  DFFPOSX1 fifo_array_reg_15__22_ ( .D(n2303), .CLK(clk), .Q(fifo_array[652])
         );
  DFFPOSX1 fifo_array_reg_15__21_ ( .D(n2302), .CLK(clk), .Q(fifo_array[651])
         );
  DFFPOSX1 fifo_array_reg_15__20_ ( .D(n2301), .CLK(clk), .Q(fifo_array[650])
         );
  DFFPOSX1 fifo_array_reg_15__19_ ( .D(n2300), .CLK(clk), .Q(fifo_array[649])
         );
  DFFPOSX1 fifo_array_reg_15__18_ ( .D(n2299), .CLK(clk), .Q(fifo_array[648])
         );
  DFFPOSX1 fifo_array_reg_15__17_ ( .D(n2298), .CLK(clk), .Q(fifo_array[647])
         );
  DFFPOSX1 fifo_array_reg_15__16_ ( .D(n2297), .CLK(clk), .Q(fifo_array[646])
         );
  DFFPOSX1 fifo_array_reg_15__15_ ( .D(n2296), .CLK(clk), .Q(fifo_array[645])
         );
  DFFPOSX1 fifo_array_reg_15__14_ ( .D(n2295), .CLK(clk), .Q(fifo_array[644])
         );
  DFFPOSX1 fifo_array_reg_15__13_ ( .D(n2294), .CLK(clk), .Q(fifo_array[643])
         );
  DFFPOSX1 fifo_array_reg_15__12_ ( .D(n2293), .CLK(clk), .Q(fifo_array[642])
         );
  DFFPOSX1 fifo_array_reg_15__11_ ( .D(n2292), .CLK(clk), .Q(fifo_array[641])
         );
  DFFPOSX1 fifo_array_reg_15__10_ ( .D(n2291), .CLK(clk), .Q(fifo_array[640])
         );
  DFFPOSX1 fifo_array_reg_15__9_ ( .D(n2290), .CLK(clk), .Q(fifo_array[639])
         );
  DFFPOSX1 fifo_array_reg_15__8_ ( .D(n2289), .CLK(clk), .Q(fifo_array[638])
         );
  DFFPOSX1 fifo_array_reg_15__7_ ( .D(n2288), .CLK(clk), .Q(fifo_array[637])
         );
  DFFPOSX1 fifo_array_reg_15__6_ ( .D(n2287), .CLK(clk), .Q(fifo_array[636])
         );
  DFFPOSX1 fifo_array_reg_15__5_ ( .D(n2286), .CLK(clk), .Q(fifo_array[635])
         );
  DFFPOSX1 fifo_array_reg_15__4_ ( .D(n2285), .CLK(clk), .Q(fifo_array[634])
         );
  DFFPOSX1 fifo_array_reg_15__3_ ( .D(n2284), .CLK(clk), .Q(fifo_array[633])
         );
  DFFPOSX1 fifo_array_reg_15__2_ ( .D(n2283), .CLK(clk), .Q(fifo_array[632])
         );
  DFFPOSX1 fifo_array_reg_15__1_ ( .D(n2282), .CLK(clk), .Q(fifo_array[631])
         );
  DFFPOSX1 fifo_array_reg_15__0_ ( .D(n2281), .CLK(clk), .Q(fifo_array[630])
         );
  DFFPOSX1 fifo_array_reg_14__41_ ( .D(n2280), .CLK(clk), .Q(fifo_array[629])
         );
  DFFPOSX1 fifo_array_reg_14__40_ ( .D(n2279), .CLK(clk), .Q(fifo_array[628])
         );
  DFFPOSX1 fifo_array_reg_14__39_ ( .D(n2278), .CLK(clk), .Q(fifo_array[627])
         );
  DFFPOSX1 fifo_array_reg_14__38_ ( .D(n2277), .CLK(clk), .Q(fifo_array[626])
         );
  DFFPOSX1 fifo_array_reg_14__37_ ( .D(n2276), .CLK(clk), .Q(fifo_array[625])
         );
  DFFPOSX1 fifo_array_reg_14__36_ ( .D(n2275), .CLK(clk), .Q(fifo_array[624])
         );
  DFFPOSX1 fifo_array_reg_14__35_ ( .D(n2274), .CLK(clk), .Q(fifo_array[623])
         );
  DFFPOSX1 fifo_array_reg_14__34_ ( .D(n2273), .CLK(clk), .Q(fifo_array[622])
         );
  DFFPOSX1 fifo_array_reg_14__33_ ( .D(n2272), .CLK(clk), .Q(fifo_array[621])
         );
  DFFPOSX1 fifo_array_reg_14__32_ ( .D(n2271), .CLK(clk), .Q(fifo_array[620])
         );
  DFFPOSX1 fifo_array_reg_14__31_ ( .D(n2270), .CLK(clk), .Q(fifo_array[619])
         );
  DFFPOSX1 fifo_array_reg_14__30_ ( .D(n2269), .CLK(clk), .Q(fifo_array[618])
         );
  DFFPOSX1 fifo_array_reg_14__29_ ( .D(n2268), .CLK(clk), .Q(fifo_array[617])
         );
  DFFPOSX1 fifo_array_reg_14__28_ ( .D(n2267), .CLK(clk), .Q(fifo_array[616])
         );
  DFFPOSX1 fifo_array_reg_14__27_ ( .D(n2266), .CLK(clk), .Q(fifo_array[615])
         );
  DFFPOSX1 fifo_array_reg_14__26_ ( .D(n2265), .CLK(clk), .Q(fifo_array[614])
         );
  DFFPOSX1 fifo_array_reg_14__25_ ( .D(n2264), .CLK(clk), .Q(fifo_array[613])
         );
  DFFPOSX1 fifo_array_reg_14__24_ ( .D(n2263), .CLK(clk), .Q(fifo_array[612])
         );
  DFFPOSX1 fifo_array_reg_14__23_ ( .D(n2262), .CLK(clk), .Q(fifo_array[611])
         );
  DFFPOSX1 fifo_array_reg_14__22_ ( .D(n2261), .CLK(clk), .Q(fifo_array[610])
         );
  DFFPOSX1 fifo_array_reg_14__21_ ( .D(n2260), .CLK(clk), .Q(fifo_array[609])
         );
  DFFPOSX1 fifo_array_reg_14__20_ ( .D(n2259), .CLK(clk), .Q(fifo_array[608])
         );
  DFFPOSX1 fifo_array_reg_14__19_ ( .D(n2258), .CLK(clk), .Q(fifo_array[607])
         );
  DFFPOSX1 fifo_array_reg_14__18_ ( .D(n2257), .CLK(clk), .Q(fifo_array[606])
         );
  DFFPOSX1 fifo_array_reg_14__17_ ( .D(n2256), .CLK(clk), .Q(fifo_array[605])
         );
  DFFPOSX1 fifo_array_reg_14__16_ ( .D(n2255), .CLK(clk), .Q(fifo_array[604])
         );
  DFFPOSX1 fifo_array_reg_14__15_ ( .D(n2254), .CLK(clk), .Q(fifo_array[603])
         );
  DFFPOSX1 fifo_array_reg_14__14_ ( .D(n2253), .CLK(clk), .Q(fifo_array[602])
         );
  DFFPOSX1 fifo_array_reg_14__13_ ( .D(n2252), .CLK(clk), .Q(fifo_array[601])
         );
  DFFPOSX1 fifo_array_reg_14__12_ ( .D(n2251), .CLK(clk), .Q(fifo_array[600])
         );
  DFFPOSX1 fifo_array_reg_14__11_ ( .D(n2250), .CLK(clk), .Q(fifo_array[599])
         );
  DFFPOSX1 fifo_array_reg_14__10_ ( .D(n2249), .CLK(clk), .Q(fifo_array[598])
         );
  DFFPOSX1 fifo_array_reg_14__9_ ( .D(n2248), .CLK(clk), .Q(fifo_array[597])
         );
  DFFPOSX1 fifo_array_reg_14__8_ ( .D(n2247), .CLK(clk), .Q(fifo_array[596])
         );
  DFFPOSX1 fifo_array_reg_14__7_ ( .D(n2246), .CLK(clk), .Q(fifo_array[595])
         );
  DFFPOSX1 fifo_array_reg_14__6_ ( .D(n2245), .CLK(clk), .Q(fifo_array[594])
         );
  DFFPOSX1 fifo_array_reg_14__5_ ( .D(n2244), .CLK(clk), .Q(fifo_array[593])
         );
  DFFPOSX1 fifo_array_reg_14__4_ ( .D(n2243), .CLK(clk), .Q(fifo_array[592])
         );
  DFFPOSX1 fifo_array_reg_14__3_ ( .D(n2242), .CLK(clk), .Q(fifo_array[591])
         );
  DFFPOSX1 fifo_array_reg_14__2_ ( .D(n2241), .CLK(clk), .Q(fifo_array[590])
         );
  DFFPOSX1 fifo_array_reg_14__1_ ( .D(n2240), .CLK(clk), .Q(fifo_array[589])
         );
  DFFPOSX1 fifo_array_reg_14__0_ ( .D(n2239), .CLK(clk), .Q(fifo_array[588])
         );
  DFFPOSX1 fifo_array_reg_13__41_ ( .D(n2238), .CLK(clk), .Q(fifo_array[587])
         );
  DFFPOSX1 fifo_array_reg_13__40_ ( .D(n2237), .CLK(clk), .Q(fifo_array[586])
         );
  DFFPOSX1 fifo_array_reg_13__39_ ( .D(n2236), .CLK(clk), .Q(fifo_array[585])
         );
  DFFPOSX1 fifo_array_reg_13__38_ ( .D(n2235), .CLK(clk), .Q(fifo_array[584])
         );
  DFFPOSX1 fifo_array_reg_13__37_ ( .D(n2234), .CLK(clk), .Q(fifo_array[583])
         );
  DFFPOSX1 fifo_array_reg_13__36_ ( .D(n2233), .CLK(clk), .Q(fifo_array[582])
         );
  DFFPOSX1 fifo_array_reg_13__35_ ( .D(n2232), .CLK(clk), .Q(fifo_array[581])
         );
  DFFPOSX1 fifo_array_reg_13__34_ ( .D(n2231), .CLK(clk), .Q(fifo_array[580])
         );
  DFFPOSX1 fifo_array_reg_13__33_ ( .D(n2230), .CLK(clk), .Q(fifo_array[579])
         );
  DFFPOSX1 fifo_array_reg_13__32_ ( .D(n2229), .CLK(clk), .Q(fifo_array[578])
         );
  DFFPOSX1 fifo_array_reg_13__31_ ( .D(n2228), .CLK(clk), .Q(fifo_array[577])
         );
  DFFPOSX1 fifo_array_reg_13__30_ ( .D(n2227), .CLK(clk), .Q(fifo_array[576])
         );
  DFFPOSX1 fifo_array_reg_13__29_ ( .D(n2226), .CLK(clk), .Q(fifo_array[575])
         );
  DFFPOSX1 fifo_array_reg_13__28_ ( .D(n2225), .CLK(clk), .Q(fifo_array[574])
         );
  DFFPOSX1 fifo_array_reg_13__27_ ( .D(n2224), .CLK(clk), .Q(fifo_array[573])
         );
  DFFPOSX1 fifo_array_reg_13__26_ ( .D(n2223), .CLK(clk), .Q(fifo_array[572])
         );
  DFFPOSX1 fifo_array_reg_13__25_ ( .D(n2222), .CLK(clk), .Q(fifo_array[571])
         );
  DFFPOSX1 fifo_array_reg_13__24_ ( .D(n2221), .CLK(clk), .Q(fifo_array[570])
         );
  DFFPOSX1 fifo_array_reg_13__23_ ( .D(n2220), .CLK(clk), .Q(fifo_array[569])
         );
  DFFPOSX1 fifo_array_reg_13__22_ ( .D(n2219), .CLK(clk), .Q(fifo_array[568])
         );
  DFFPOSX1 fifo_array_reg_13__21_ ( .D(n2218), .CLK(clk), .Q(fifo_array[567])
         );
  DFFPOSX1 fifo_array_reg_13__20_ ( .D(n2217), .CLK(clk), .Q(fifo_array[566])
         );
  DFFPOSX1 fifo_array_reg_13__19_ ( .D(n2216), .CLK(clk), .Q(fifo_array[565])
         );
  DFFPOSX1 fifo_array_reg_13__18_ ( .D(n2215), .CLK(clk), .Q(fifo_array[564])
         );
  DFFPOSX1 fifo_array_reg_13__17_ ( .D(n2214), .CLK(clk), .Q(fifo_array[563])
         );
  DFFPOSX1 fifo_array_reg_13__16_ ( .D(n2213), .CLK(clk), .Q(fifo_array[562])
         );
  DFFPOSX1 fifo_array_reg_13__15_ ( .D(n2212), .CLK(clk), .Q(fifo_array[561])
         );
  DFFPOSX1 fifo_array_reg_13__14_ ( .D(n2211), .CLK(clk), .Q(fifo_array[560])
         );
  DFFPOSX1 fifo_array_reg_13__13_ ( .D(n2210), .CLK(clk), .Q(fifo_array[559])
         );
  DFFPOSX1 fifo_array_reg_13__12_ ( .D(n2209), .CLK(clk), .Q(fifo_array[558])
         );
  DFFPOSX1 fifo_array_reg_13__11_ ( .D(n2208), .CLK(clk), .Q(fifo_array[557])
         );
  DFFPOSX1 fifo_array_reg_13__10_ ( .D(n2207), .CLK(clk), .Q(fifo_array[556])
         );
  DFFPOSX1 fifo_array_reg_13__9_ ( .D(n2206), .CLK(clk), .Q(fifo_array[555])
         );
  DFFPOSX1 fifo_array_reg_13__8_ ( .D(n2205), .CLK(clk), .Q(fifo_array[554])
         );
  DFFPOSX1 fifo_array_reg_13__7_ ( .D(n2204), .CLK(clk), .Q(fifo_array[553])
         );
  DFFPOSX1 fifo_array_reg_13__6_ ( .D(n2203), .CLK(clk), .Q(fifo_array[552])
         );
  DFFPOSX1 fifo_array_reg_13__5_ ( .D(n2202), .CLK(clk), .Q(fifo_array[551])
         );
  DFFPOSX1 fifo_array_reg_13__4_ ( .D(n2201), .CLK(clk), .Q(fifo_array[550])
         );
  DFFPOSX1 fifo_array_reg_13__3_ ( .D(n2200), .CLK(clk), .Q(fifo_array[549])
         );
  DFFPOSX1 fifo_array_reg_13__2_ ( .D(n2199), .CLK(clk), .Q(fifo_array[548])
         );
  DFFPOSX1 fifo_array_reg_13__1_ ( .D(n2198), .CLK(clk), .Q(fifo_array[547])
         );
  DFFPOSX1 fifo_array_reg_13__0_ ( .D(n2197), .CLK(clk), .Q(fifo_array[546])
         );
  DFFPOSX1 fifo_array_reg_12__41_ ( .D(n2196), .CLK(clk), .Q(fifo_array[545])
         );
  DFFPOSX1 fifo_array_reg_12__40_ ( .D(n2195), .CLK(clk), .Q(fifo_array[544])
         );
  DFFPOSX1 fifo_array_reg_12__39_ ( .D(n2194), .CLK(clk), .Q(fifo_array[543])
         );
  DFFPOSX1 fifo_array_reg_12__38_ ( .D(n2193), .CLK(clk), .Q(fifo_array[542])
         );
  DFFPOSX1 fifo_array_reg_12__37_ ( .D(n2192), .CLK(clk), .Q(fifo_array[541])
         );
  DFFPOSX1 fifo_array_reg_12__36_ ( .D(n2191), .CLK(clk), .Q(fifo_array[540])
         );
  DFFPOSX1 fifo_array_reg_12__35_ ( .D(n2190), .CLK(clk), .Q(fifo_array[539])
         );
  DFFPOSX1 fifo_array_reg_12__34_ ( .D(n2189), .CLK(clk), .Q(fifo_array[538])
         );
  DFFPOSX1 fifo_array_reg_12__33_ ( .D(n2188), .CLK(clk), .Q(fifo_array[537])
         );
  DFFPOSX1 fifo_array_reg_12__32_ ( .D(n2187), .CLK(clk), .Q(fifo_array[536])
         );
  DFFPOSX1 fifo_array_reg_12__31_ ( .D(n2186), .CLK(clk), .Q(fifo_array[535])
         );
  DFFPOSX1 fifo_array_reg_12__30_ ( .D(n2185), .CLK(clk), .Q(fifo_array[534])
         );
  DFFPOSX1 fifo_array_reg_12__29_ ( .D(n2184), .CLK(clk), .Q(fifo_array[533])
         );
  DFFPOSX1 fifo_array_reg_12__28_ ( .D(n2183), .CLK(clk), .Q(fifo_array[532])
         );
  DFFPOSX1 fifo_array_reg_12__27_ ( .D(n2182), .CLK(clk), .Q(fifo_array[531])
         );
  DFFPOSX1 fifo_array_reg_12__26_ ( .D(n2181), .CLK(clk), .Q(fifo_array[530])
         );
  DFFPOSX1 fifo_array_reg_12__25_ ( .D(n2180), .CLK(clk), .Q(fifo_array[529])
         );
  DFFPOSX1 fifo_array_reg_12__24_ ( .D(n2179), .CLK(clk), .Q(fifo_array[528])
         );
  DFFPOSX1 fifo_array_reg_12__23_ ( .D(n2178), .CLK(clk), .Q(fifo_array[527])
         );
  DFFPOSX1 fifo_array_reg_12__22_ ( .D(n2177), .CLK(clk), .Q(fifo_array[526])
         );
  DFFPOSX1 fifo_array_reg_12__21_ ( .D(n2176), .CLK(clk), .Q(fifo_array[525])
         );
  DFFPOSX1 fifo_array_reg_12__20_ ( .D(n2175), .CLK(clk), .Q(fifo_array[524])
         );
  DFFPOSX1 fifo_array_reg_12__19_ ( .D(n2174), .CLK(clk), .Q(fifo_array[523])
         );
  DFFPOSX1 fifo_array_reg_12__18_ ( .D(n2173), .CLK(clk), .Q(fifo_array[522])
         );
  DFFPOSX1 fifo_array_reg_12__17_ ( .D(n2172), .CLK(clk), .Q(fifo_array[521])
         );
  DFFPOSX1 fifo_array_reg_12__16_ ( .D(n2171), .CLK(clk), .Q(fifo_array[520])
         );
  DFFPOSX1 fifo_array_reg_12__15_ ( .D(n2170), .CLK(clk), .Q(fifo_array[519])
         );
  DFFPOSX1 fifo_array_reg_12__14_ ( .D(n2169), .CLK(clk), .Q(fifo_array[518])
         );
  DFFPOSX1 fifo_array_reg_12__13_ ( .D(n2168), .CLK(clk), .Q(fifo_array[517])
         );
  DFFPOSX1 fifo_array_reg_12__12_ ( .D(n2167), .CLK(clk), .Q(fifo_array[516])
         );
  DFFPOSX1 fifo_array_reg_12__11_ ( .D(n2166), .CLK(clk), .Q(fifo_array[515])
         );
  DFFPOSX1 fifo_array_reg_12__10_ ( .D(n2165), .CLK(clk), .Q(fifo_array[514])
         );
  DFFPOSX1 fifo_array_reg_12__9_ ( .D(n2164), .CLK(clk), .Q(fifo_array[513])
         );
  DFFPOSX1 fifo_array_reg_12__8_ ( .D(n2163), .CLK(clk), .Q(fifo_array[512])
         );
  DFFPOSX1 fifo_array_reg_12__7_ ( .D(n2162), .CLK(clk), .Q(fifo_array[511])
         );
  DFFPOSX1 fifo_array_reg_12__6_ ( .D(n2161), .CLK(clk), .Q(fifo_array[510])
         );
  DFFPOSX1 fifo_array_reg_12__5_ ( .D(n2160), .CLK(clk), .Q(fifo_array[509])
         );
  DFFPOSX1 fifo_array_reg_12__4_ ( .D(n2159), .CLK(clk), .Q(fifo_array[508])
         );
  DFFPOSX1 fifo_array_reg_12__3_ ( .D(n2158), .CLK(clk), .Q(fifo_array[507])
         );
  DFFPOSX1 fifo_array_reg_12__2_ ( .D(n2157), .CLK(clk), .Q(fifo_array[506])
         );
  DFFPOSX1 fifo_array_reg_12__1_ ( .D(n2156), .CLK(clk), .Q(fifo_array[505])
         );
  DFFPOSX1 fifo_array_reg_12__0_ ( .D(n2155), .CLK(clk), .Q(fifo_array[504])
         );
  DFFPOSX1 fifo_array_reg_11__41_ ( .D(n2154), .CLK(clk), .Q(fifo_array[503])
         );
  DFFPOSX1 fifo_array_reg_11__40_ ( .D(n2153), .CLK(clk), .Q(fifo_array[502])
         );
  DFFPOSX1 fifo_array_reg_11__39_ ( .D(n2152), .CLK(clk), .Q(fifo_array[501])
         );
  DFFPOSX1 fifo_array_reg_11__38_ ( .D(n2151), .CLK(clk), .Q(fifo_array[500])
         );
  DFFPOSX1 fifo_array_reg_11__37_ ( .D(n2150), .CLK(clk), .Q(fifo_array[499])
         );
  DFFPOSX1 fifo_array_reg_11__36_ ( .D(n2149), .CLK(clk), .Q(fifo_array[498])
         );
  DFFPOSX1 fifo_array_reg_11__35_ ( .D(n2148), .CLK(clk), .Q(fifo_array[497])
         );
  DFFPOSX1 fifo_array_reg_11__34_ ( .D(n2147), .CLK(clk), .Q(fifo_array[496])
         );
  DFFPOSX1 fifo_array_reg_11__33_ ( .D(n2146), .CLK(clk), .Q(fifo_array[495])
         );
  DFFPOSX1 fifo_array_reg_11__32_ ( .D(n2145), .CLK(clk), .Q(fifo_array[494])
         );
  DFFPOSX1 fifo_array_reg_11__31_ ( .D(n2144), .CLK(clk), .Q(fifo_array[493])
         );
  DFFPOSX1 fifo_array_reg_11__30_ ( .D(n2143), .CLK(clk), .Q(fifo_array[492])
         );
  DFFPOSX1 fifo_array_reg_11__29_ ( .D(n2142), .CLK(clk), .Q(fifo_array[491])
         );
  DFFPOSX1 fifo_array_reg_11__28_ ( .D(n2141), .CLK(clk), .Q(fifo_array[490])
         );
  DFFPOSX1 fifo_array_reg_11__27_ ( .D(n2140), .CLK(clk), .Q(fifo_array[489])
         );
  DFFPOSX1 fifo_array_reg_11__26_ ( .D(n2139), .CLK(clk), .Q(fifo_array[488])
         );
  DFFPOSX1 fifo_array_reg_11__25_ ( .D(n2138), .CLK(clk), .Q(fifo_array[487])
         );
  DFFPOSX1 fifo_array_reg_11__24_ ( .D(n2137), .CLK(clk), .Q(fifo_array[486])
         );
  DFFPOSX1 fifo_array_reg_11__23_ ( .D(n2136), .CLK(clk), .Q(fifo_array[485])
         );
  DFFPOSX1 fifo_array_reg_11__22_ ( .D(n2135), .CLK(clk), .Q(fifo_array[484])
         );
  DFFPOSX1 fifo_array_reg_11__21_ ( .D(n2134), .CLK(clk), .Q(fifo_array[483])
         );
  DFFPOSX1 fifo_array_reg_11__20_ ( .D(n2133), .CLK(clk), .Q(fifo_array[482])
         );
  DFFPOSX1 fifo_array_reg_11__19_ ( .D(n2132), .CLK(clk), .Q(fifo_array[481])
         );
  DFFPOSX1 fifo_array_reg_11__18_ ( .D(n2131), .CLK(clk), .Q(fifo_array[480])
         );
  DFFPOSX1 fifo_array_reg_11__17_ ( .D(n2130), .CLK(clk), .Q(fifo_array[479])
         );
  DFFPOSX1 fifo_array_reg_11__16_ ( .D(n2129), .CLK(clk), .Q(fifo_array[478])
         );
  DFFPOSX1 fifo_array_reg_11__15_ ( .D(n2128), .CLK(clk), .Q(fifo_array[477])
         );
  DFFPOSX1 fifo_array_reg_11__14_ ( .D(n2127), .CLK(clk), .Q(fifo_array[476])
         );
  DFFPOSX1 fifo_array_reg_11__13_ ( .D(n2126), .CLK(clk), .Q(fifo_array[475])
         );
  DFFPOSX1 fifo_array_reg_11__12_ ( .D(n2125), .CLK(clk), .Q(fifo_array[474])
         );
  DFFPOSX1 fifo_array_reg_11__11_ ( .D(n2124), .CLK(clk), .Q(fifo_array[473])
         );
  DFFPOSX1 fifo_array_reg_11__10_ ( .D(n2123), .CLK(clk), .Q(fifo_array[472])
         );
  DFFPOSX1 fifo_array_reg_11__9_ ( .D(n2122), .CLK(clk), .Q(fifo_array[471])
         );
  DFFPOSX1 fifo_array_reg_11__8_ ( .D(n2121), .CLK(clk), .Q(fifo_array[470])
         );
  DFFPOSX1 fifo_array_reg_11__7_ ( .D(n2120), .CLK(clk), .Q(fifo_array[469])
         );
  DFFPOSX1 fifo_array_reg_11__6_ ( .D(n2119), .CLK(clk), .Q(fifo_array[468])
         );
  DFFPOSX1 fifo_array_reg_11__5_ ( .D(n2118), .CLK(clk), .Q(fifo_array[467])
         );
  DFFPOSX1 fifo_array_reg_11__4_ ( .D(n2117), .CLK(clk), .Q(fifo_array[466])
         );
  DFFPOSX1 fifo_array_reg_11__3_ ( .D(n2116), .CLK(clk), .Q(fifo_array[465])
         );
  DFFPOSX1 fifo_array_reg_11__2_ ( .D(n2115), .CLK(clk), .Q(fifo_array[464])
         );
  DFFPOSX1 fifo_array_reg_11__1_ ( .D(n2114), .CLK(clk), .Q(fifo_array[463])
         );
  DFFPOSX1 fifo_array_reg_11__0_ ( .D(n2113), .CLK(clk), .Q(fifo_array[462])
         );
  DFFPOSX1 fifo_array_reg_10__41_ ( .D(n2112), .CLK(clk), .Q(fifo_array[461])
         );
  DFFPOSX1 fifo_array_reg_10__40_ ( .D(n2111), .CLK(clk), .Q(fifo_array[460])
         );
  DFFPOSX1 fifo_array_reg_10__39_ ( .D(n2110), .CLK(clk), .Q(fifo_array[459])
         );
  DFFPOSX1 fifo_array_reg_10__38_ ( .D(n2109), .CLK(clk), .Q(fifo_array[458])
         );
  DFFPOSX1 fifo_array_reg_10__37_ ( .D(n2108), .CLK(clk), .Q(fifo_array[457])
         );
  DFFPOSX1 fifo_array_reg_10__36_ ( .D(n2107), .CLK(clk), .Q(fifo_array[456])
         );
  DFFPOSX1 fifo_array_reg_10__35_ ( .D(n2106), .CLK(clk), .Q(fifo_array[455])
         );
  DFFPOSX1 fifo_array_reg_10__34_ ( .D(n2105), .CLK(clk), .Q(fifo_array[454])
         );
  DFFPOSX1 fifo_array_reg_10__33_ ( .D(n2104), .CLK(clk), .Q(fifo_array[453])
         );
  DFFPOSX1 fifo_array_reg_10__32_ ( .D(n2103), .CLK(clk), .Q(fifo_array[452])
         );
  DFFPOSX1 fifo_array_reg_10__31_ ( .D(n2102), .CLK(clk), .Q(fifo_array[451])
         );
  DFFPOSX1 fifo_array_reg_10__30_ ( .D(n2101), .CLK(clk), .Q(fifo_array[450])
         );
  DFFPOSX1 fifo_array_reg_10__29_ ( .D(n2100), .CLK(clk), .Q(fifo_array[449])
         );
  DFFPOSX1 fifo_array_reg_10__28_ ( .D(n2099), .CLK(clk), .Q(fifo_array[448])
         );
  DFFPOSX1 fifo_array_reg_10__27_ ( .D(n2098), .CLK(clk), .Q(fifo_array[447])
         );
  DFFPOSX1 fifo_array_reg_10__26_ ( .D(n2097), .CLK(clk), .Q(fifo_array[446])
         );
  DFFPOSX1 fifo_array_reg_10__25_ ( .D(n2096), .CLK(clk), .Q(fifo_array[445])
         );
  DFFPOSX1 fifo_array_reg_10__24_ ( .D(n2095), .CLK(clk), .Q(fifo_array[444])
         );
  DFFPOSX1 fifo_array_reg_10__23_ ( .D(n2094), .CLK(clk), .Q(fifo_array[443])
         );
  DFFPOSX1 fifo_array_reg_10__22_ ( .D(n2093), .CLK(clk), .Q(fifo_array[442])
         );
  DFFPOSX1 fifo_array_reg_10__21_ ( .D(n2092), .CLK(clk), .Q(fifo_array[441])
         );
  DFFPOSX1 fifo_array_reg_10__20_ ( .D(n2091), .CLK(clk), .Q(fifo_array[440])
         );
  DFFPOSX1 fifo_array_reg_10__19_ ( .D(n2090), .CLK(clk), .Q(fifo_array[439])
         );
  DFFPOSX1 fifo_array_reg_10__18_ ( .D(n2089), .CLK(clk), .Q(fifo_array[438])
         );
  DFFPOSX1 fifo_array_reg_10__17_ ( .D(n2088), .CLK(clk), .Q(fifo_array[437])
         );
  DFFPOSX1 fifo_array_reg_10__16_ ( .D(n2087), .CLK(clk), .Q(fifo_array[436])
         );
  DFFPOSX1 fifo_array_reg_10__15_ ( .D(n2086), .CLK(clk), .Q(fifo_array[435])
         );
  DFFPOSX1 fifo_array_reg_10__14_ ( .D(n2085), .CLK(clk), .Q(fifo_array[434])
         );
  DFFPOSX1 fifo_array_reg_10__13_ ( .D(n2084), .CLK(clk), .Q(fifo_array[433])
         );
  DFFPOSX1 fifo_array_reg_10__12_ ( .D(n2083), .CLK(clk), .Q(fifo_array[432])
         );
  DFFPOSX1 fifo_array_reg_10__11_ ( .D(n2082), .CLK(clk), .Q(fifo_array[431])
         );
  DFFPOSX1 fifo_array_reg_10__10_ ( .D(n2081), .CLK(clk), .Q(fifo_array[430])
         );
  DFFPOSX1 fifo_array_reg_10__9_ ( .D(n2080), .CLK(clk), .Q(fifo_array[429])
         );
  DFFPOSX1 fifo_array_reg_10__8_ ( .D(n2079), .CLK(clk), .Q(fifo_array[428])
         );
  DFFPOSX1 fifo_array_reg_10__7_ ( .D(n2078), .CLK(clk), .Q(fifo_array[427])
         );
  DFFPOSX1 fifo_array_reg_10__6_ ( .D(n2077), .CLK(clk), .Q(fifo_array[426])
         );
  DFFPOSX1 fifo_array_reg_10__5_ ( .D(n2076), .CLK(clk), .Q(fifo_array[425])
         );
  DFFPOSX1 fifo_array_reg_10__4_ ( .D(n2075), .CLK(clk), .Q(fifo_array[424])
         );
  DFFPOSX1 fifo_array_reg_10__3_ ( .D(n2074), .CLK(clk), .Q(fifo_array[423])
         );
  DFFPOSX1 fifo_array_reg_10__2_ ( .D(n2073), .CLK(clk), .Q(fifo_array[422])
         );
  DFFPOSX1 fifo_array_reg_10__1_ ( .D(n2072), .CLK(clk), .Q(fifo_array[421])
         );
  DFFPOSX1 fifo_array_reg_10__0_ ( .D(n2071), .CLK(clk), .Q(fifo_array[420])
         );
  DFFPOSX1 fifo_array_reg_9__41_ ( .D(n2070), .CLK(clk), .Q(fifo_array[419])
         );
  DFFPOSX1 fifo_array_reg_9__40_ ( .D(n2069), .CLK(clk), .Q(fifo_array[418])
         );
  DFFPOSX1 fifo_array_reg_9__39_ ( .D(n2068), .CLK(clk), .Q(fifo_array[417])
         );
  DFFPOSX1 fifo_array_reg_9__38_ ( .D(n2067), .CLK(clk), .Q(fifo_array[416])
         );
  DFFPOSX1 fifo_array_reg_9__37_ ( .D(n2066), .CLK(clk), .Q(fifo_array[415])
         );
  DFFPOSX1 fifo_array_reg_9__36_ ( .D(n2065), .CLK(clk), .Q(fifo_array[414])
         );
  DFFPOSX1 fifo_array_reg_9__35_ ( .D(n2064), .CLK(clk), .Q(fifo_array[413])
         );
  DFFPOSX1 fifo_array_reg_9__34_ ( .D(n2063), .CLK(clk), .Q(fifo_array[412])
         );
  DFFPOSX1 fifo_array_reg_9__33_ ( .D(n2062), .CLK(clk), .Q(fifo_array[411])
         );
  DFFPOSX1 fifo_array_reg_9__32_ ( .D(n2061), .CLK(clk), .Q(fifo_array[410])
         );
  DFFPOSX1 fifo_array_reg_9__31_ ( .D(n2060), .CLK(clk), .Q(fifo_array[409])
         );
  DFFPOSX1 fifo_array_reg_9__30_ ( .D(n2059), .CLK(clk), .Q(fifo_array[408])
         );
  DFFPOSX1 fifo_array_reg_9__29_ ( .D(n2058), .CLK(clk), .Q(fifo_array[407])
         );
  DFFPOSX1 fifo_array_reg_9__28_ ( .D(n2057), .CLK(clk), .Q(fifo_array[406])
         );
  DFFPOSX1 fifo_array_reg_9__27_ ( .D(n2056), .CLK(clk), .Q(fifo_array[405])
         );
  DFFPOSX1 fifo_array_reg_9__26_ ( .D(n2055), .CLK(clk), .Q(fifo_array[404])
         );
  DFFPOSX1 fifo_array_reg_9__25_ ( .D(n2054), .CLK(clk), .Q(fifo_array[403])
         );
  DFFPOSX1 fifo_array_reg_9__24_ ( .D(n2053), .CLK(clk), .Q(fifo_array[402])
         );
  DFFPOSX1 fifo_array_reg_9__23_ ( .D(n2052), .CLK(clk), .Q(fifo_array[401])
         );
  DFFPOSX1 fifo_array_reg_9__22_ ( .D(n2051), .CLK(clk), .Q(fifo_array[400])
         );
  DFFPOSX1 fifo_array_reg_9__21_ ( .D(n2050), .CLK(clk), .Q(fifo_array[399])
         );
  DFFPOSX1 fifo_array_reg_9__20_ ( .D(n2049), .CLK(clk), .Q(fifo_array[398])
         );
  DFFPOSX1 fifo_array_reg_9__19_ ( .D(n2048), .CLK(clk), .Q(fifo_array[397])
         );
  DFFPOSX1 fifo_array_reg_9__18_ ( .D(n2047), .CLK(clk), .Q(fifo_array[396])
         );
  DFFPOSX1 fifo_array_reg_9__17_ ( .D(n2046), .CLK(clk), .Q(fifo_array[395])
         );
  DFFPOSX1 fifo_array_reg_9__16_ ( .D(n2045), .CLK(clk), .Q(fifo_array[394])
         );
  DFFPOSX1 fifo_array_reg_9__15_ ( .D(n2044), .CLK(clk), .Q(fifo_array[393])
         );
  DFFPOSX1 fifo_array_reg_9__14_ ( .D(n2043), .CLK(clk), .Q(fifo_array[392])
         );
  DFFPOSX1 fifo_array_reg_9__13_ ( .D(n2042), .CLK(clk), .Q(fifo_array[391])
         );
  DFFPOSX1 fifo_array_reg_9__12_ ( .D(n2041), .CLK(clk), .Q(fifo_array[390])
         );
  DFFPOSX1 fifo_array_reg_9__11_ ( .D(n2040), .CLK(clk), .Q(fifo_array[389])
         );
  DFFPOSX1 fifo_array_reg_9__10_ ( .D(n2039), .CLK(clk), .Q(fifo_array[388])
         );
  DFFPOSX1 fifo_array_reg_9__9_ ( .D(n2038), .CLK(clk), .Q(fifo_array[387]) );
  DFFPOSX1 fifo_array_reg_9__8_ ( .D(n2037), .CLK(clk), .Q(fifo_array[386]) );
  DFFPOSX1 fifo_array_reg_9__7_ ( .D(n2036), .CLK(clk), .Q(fifo_array[385]) );
  DFFPOSX1 fifo_array_reg_9__6_ ( .D(n2035), .CLK(clk), .Q(fifo_array[384]) );
  DFFPOSX1 fifo_array_reg_9__5_ ( .D(n2034), .CLK(clk), .Q(fifo_array[383]) );
  DFFPOSX1 fifo_array_reg_9__4_ ( .D(n2033), .CLK(clk), .Q(fifo_array[382]) );
  DFFPOSX1 fifo_array_reg_9__3_ ( .D(n2032), .CLK(clk), .Q(fifo_array[381]) );
  DFFPOSX1 fifo_array_reg_9__2_ ( .D(n2031), .CLK(clk), .Q(fifo_array[380]) );
  DFFPOSX1 fifo_array_reg_9__1_ ( .D(n2030), .CLK(clk), .Q(fifo_array[379]) );
  DFFPOSX1 fifo_array_reg_9__0_ ( .D(n2029), .CLK(clk), .Q(fifo_array[378]) );
  DFFPOSX1 fifo_array_reg_8__41_ ( .D(n2028), .CLK(clk), .Q(fifo_array[377])
         );
  DFFPOSX1 fifo_array_reg_8__40_ ( .D(n2027), .CLK(clk), .Q(fifo_array[376])
         );
  DFFPOSX1 fifo_array_reg_8__39_ ( .D(n2026), .CLK(clk), .Q(fifo_array[375])
         );
  DFFPOSX1 fifo_array_reg_8__38_ ( .D(n2025), .CLK(clk), .Q(fifo_array[374])
         );
  DFFPOSX1 fifo_array_reg_8__37_ ( .D(n2024), .CLK(clk), .Q(fifo_array[373])
         );
  DFFPOSX1 fifo_array_reg_8__36_ ( .D(n2023), .CLK(clk), .Q(fifo_array[372])
         );
  DFFPOSX1 fifo_array_reg_8__35_ ( .D(n2022), .CLK(clk), .Q(fifo_array[371])
         );
  DFFPOSX1 fifo_array_reg_8__34_ ( .D(n2021), .CLK(clk), .Q(fifo_array[370])
         );
  DFFPOSX1 fifo_array_reg_8__33_ ( .D(n2020), .CLK(clk), .Q(fifo_array[369])
         );
  DFFPOSX1 fifo_array_reg_8__32_ ( .D(n2019), .CLK(clk), .Q(fifo_array[368])
         );
  DFFPOSX1 fifo_array_reg_8__31_ ( .D(n2018), .CLK(clk), .Q(fifo_array[367])
         );
  DFFPOSX1 fifo_array_reg_8__30_ ( .D(n2017), .CLK(clk), .Q(fifo_array[366])
         );
  DFFPOSX1 fifo_array_reg_8__29_ ( .D(n2016), .CLK(clk), .Q(fifo_array[365])
         );
  DFFPOSX1 fifo_array_reg_8__28_ ( .D(n2015), .CLK(clk), .Q(fifo_array[364])
         );
  DFFPOSX1 fifo_array_reg_8__27_ ( .D(n2014), .CLK(clk), .Q(fifo_array[363])
         );
  DFFPOSX1 fifo_array_reg_8__26_ ( .D(n2013), .CLK(clk), .Q(fifo_array[362])
         );
  DFFPOSX1 fifo_array_reg_8__25_ ( .D(n2012), .CLK(clk), .Q(fifo_array[361])
         );
  DFFPOSX1 fifo_array_reg_8__24_ ( .D(n2011), .CLK(clk), .Q(fifo_array[360])
         );
  DFFPOSX1 fifo_array_reg_8__23_ ( .D(n2010), .CLK(clk), .Q(fifo_array[359])
         );
  DFFPOSX1 fifo_array_reg_8__22_ ( .D(n2009), .CLK(clk), .Q(fifo_array[358])
         );
  DFFPOSX1 fifo_array_reg_8__21_ ( .D(n2008), .CLK(clk), .Q(fifo_array[357])
         );
  DFFPOSX1 fifo_array_reg_8__20_ ( .D(n2007), .CLK(clk), .Q(fifo_array[356])
         );
  DFFPOSX1 fifo_array_reg_8__19_ ( .D(n2006), .CLK(clk), .Q(fifo_array[355])
         );
  DFFPOSX1 fifo_array_reg_8__18_ ( .D(n2005), .CLK(clk), .Q(fifo_array[354])
         );
  DFFPOSX1 fifo_array_reg_8__17_ ( .D(n2004), .CLK(clk), .Q(fifo_array[353])
         );
  DFFPOSX1 fifo_array_reg_8__16_ ( .D(n2003), .CLK(clk), .Q(fifo_array[352])
         );
  DFFPOSX1 fifo_array_reg_8__15_ ( .D(n2002), .CLK(clk), .Q(fifo_array[351])
         );
  DFFPOSX1 fifo_array_reg_8__14_ ( .D(n2001), .CLK(clk), .Q(fifo_array[350])
         );
  DFFPOSX1 fifo_array_reg_8__13_ ( .D(n2000), .CLK(clk), .Q(fifo_array[349])
         );
  DFFPOSX1 fifo_array_reg_8__12_ ( .D(n1999), .CLK(clk), .Q(fifo_array[348])
         );
  DFFPOSX1 fifo_array_reg_8__11_ ( .D(n1998), .CLK(clk), .Q(fifo_array[347])
         );
  DFFPOSX1 fifo_array_reg_8__10_ ( .D(n1997), .CLK(clk), .Q(fifo_array[346])
         );
  DFFPOSX1 fifo_array_reg_8__9_ ( .D(n1996), .CLK(clk), .Q(fifo_array[345]) );
  DFFPOSX1 fifo_array_reg_8__8_ ( .D(n1995), .CLK(clk), .Q(fifo_array[344]) );
  DFFPOSX1 fifo_array_reg_8__7_ ( .D(n1994), .CLK(clk), .Q(fifo_array[343]) );
  DFFPOSX1 fifo_array_reg_8__6_ ( .D(n1993), .CLK(clk), .Q(fifo_array[342]) );
  DFFPOSX1 fifo_array_reg_8__5_ ( .D(n1992), .CLK(clk), .Q(fifo_array[341]) );
  DFFPOSX1 fifo_array_reg_8__4_ ( .D(n1991), .CLK(clk), .Q(fifo_array[340]) );
  DFFPOSX1 fifo_array_reg_8__3_ ( .D(n1990), .CLK(clk), .Q(fifo_array[339]) );
  DFFPOSX1 fifo_array_reg_8__2_ ( .D(n1989), .CLK(clk), .Q(fifo_array[338]) );
  DFFPOSX1 fifo_array_reg_8__1_ ( .D(n1988), .CLK(clk), .Q(fifo_array[337]) );
  DFFPOSX1 fifo_array_reg_8__0_ ( .D(n1987), .CLK(clk), .Q(fifo_array[336]) );
  DFFPOSX1 fifo_array_reg_7__41_ ( .D(n1986), .CLK(clk), .Q(fifo_array[335])
         );
  DFFPOSX1 fifo_array_reg_7__40_ ( .D(n1985), .CLK(clk), .Q(fifo_array[334])
         );
  DFFPOSX1 fifo_array_reg_7__39_ ( .D(n1984), .CLK(clk), .Q(fifo_array[333])
         );
  DFFPOSX1 fifo_array_reg_7__38_ ( .D(n1983), .CLK(clk), .Q(fifo_array[332])
         );
  DFFPOSX1 fifo_array_reg_7__37_ ( .D(n1982), .CLK(clk), .Q(fifo_array[331])
         );
  DFFPOSX1 fifo_array_reg_7__36_ ( .D(n1981), .CLK(clk), .Q(fifo_array[330])
         );
  DFFPOSX1 fifo_array_reg_7__35_ ( .D(n1980), .CLK(clk), .Q(fifo_array[329])
         );
  DFFPOSX1 fifo_array_reg_7__34_ ( .D(n1979), .CLK(clk), .Q(fifo_array[328])
         );
  DFFPOSX1 fifo_array_reg_7__33_ ( .D(n1978), .CLK(clk), .Q(fifo_array[327])
         );
  DFFPOSX1 fifo_array_reg_7__32_ ( .D(n1977), .CLK(clk), .Q(fifo_array[326])
         );
  DFFPOSX1 fifo_array_reg_7__31_ ( .D(n1976), .CLK(clk), .Q(fifo_array[325])
         );
  DFFPOSX1 fifo_array_reg_7__30_ ( .D(n1975), .CLK(clk), .Q(fifo_array[324])
         );
  DFFPOSX1 fifo_array_reg_7__29_ ( .D(n1974), .CLK(clk), .Q(fifo_array[323])
         );
  DFFPOSX1 fifo_array_reg_7__28_ ( .D(n1973), .CLK(clk), .Q(fifo_array[322])
         );
  DFFPOSX1 fifo_array_reg_7__27_ ( .D(n1972), .CLK(clk), .Q(fifo_array[321])
         );
  DFFPOSX1 fifo_array_reg_7__26_ ( .D(n1971), .CLK(clk), .Q(fifo_array[320])
         );
  DFFPOSX1 fifo_array_reg_7__25_ ( .D(n1970), .CLK(clk), .Q(fifo_array[319])
         );
  DFFPOSX1 fifo_array_reg_7__24_ ( .D(n1969), .CLK(clk), .Q(fifo_array[318])
         );
  DFFPOSX1 fifo_array_reg_7__23_ ( .D(n1968), .CLK(clk), .Q(fifo_array[317])
         );
  DFFPOSX1 fifo_array_reg_7__22_ ( .D(n1967), .CLK(clk), .Q(fifo_array[316])
         );
  DFFPOSX1 fifo_array_reg_7__21_ ( .D(n1966), .CLK(clk), .Q(fifo_array[315])
         );
  DFFPOSX1 fifo_array_reg_7__20_ ( .D(n1965), .CLK(clk), .Q(fifo_array[314])
         );
  DFFPOSX1 fifo_array_reg_7__19_ ( .D(n1964), .CLK(clk), .Q(fifo_array[313])
         );
  DFFPOSX1 fifo_array_reg_7__18_ ( .D(n1963), .CLK(clk), .Q(fifo_array[312])
         );
  DFFPOSX1 fifo_array_reg_7__17_ ( .D(n1962), .CLK(clk), .Q(fifo_array[311])
         );
  DFFPOSX1 fifo_array_reg_7__16_ ( .D(n1961), .CLK(clk), .Q(fifo_array[310])
         );
  DFFPOSX1 fifo_array_reg_7__15_ ( .D(n1960), .CLK(clk), .Q(fifo_array[309])
         );
  DFFPOSX1 fifo_array_reg_7__14_ ( .D(n1959), .CLK(clk), .Q(fifo_array[308])
         );
  DFFPOSX1 fifo_array_reg_7__13_ ( .D(n1958), .CLK(clk), .Q(fifo_array[307])
         );
  DFFPOSX1 fifo_array_reg_7__12_ ( .D(n1957), .CLK(clk), .Q(fifo_array[306])
         );
  DFFPOSX1 fifo_array_reg_7__11_ ( .D(n1956), .CLK(clk), .Q(fifo_array[305])
         );
  DFFPOSX1 fifo_array_reg_7__10_ ( .D(n1955), .CLK(clk), .Q(fifo_array[304])
         );
  DFFPOSX1 fifo_array_reg_7__9_ ( .D(n1954), .CLK(clk), .Q(fifo_array[303]) );
  DFFPOSX1 fifo_array_reg_7__8_ ( .D(n1953), .CLK(clk), .Q(fifo_array[302]) );
  DFFPOSX1 fifo_array_reg_7__7_ ( .D(n1952), .CLK(clk), .Q(fifo_array[301]) );
  DFFPOSX1 fifo_array_reg_7__6_ ( .D(n1951), .CLK(clk), .Q(fifo_array[300]) );
  DFFPOSX1 fifo_array_reg_7__5_ ( .D(n1950), .CLK(clk), .Q(fifo_array[299]) );
  DFFPOSX1 fifo_array_reg_7__4_ ( .D(n1949), .CLK(clk), .Q(fifo_array[298]) );
  DFFPOSX1 fifo_array_reg_7__3_ ( .D(n1948), .CLK(clk), .Q(fifo_array[297]) );
  DFFPOSX1 fifo_array_reg_7__2_ ( .D(n1947), .CLK(clk), .Q(fifo_array[296]) );
  DFFPOSX1 fifo_array_reg_7__1_ ( .D(n1946), .CLK(clk), .Q(fifo_array[295]) );
  DFFPOSX1 fifo_array_reg_7__0_ ( .D(n1945), .CLK(clk), .Q(fifo_array[294]) );
  DFFPOSX1 fifo_array_reg_6__41_ ( .D(n1944), .CLK(clk), .Q(fifo_array[293])
         );
  DFFPOSX1 fifo_array_reg_6__40_ ( .D(n1943), .CLK(clk), .Q(fifo_array[292])
         );
  DFFPOSX1 fifo_array_reg_6__39_ ( .D(n1942), .CLK(clk), .Q(fifo_array[291])
         );
  DFFPOSX1 fifo_array_reg_6__38_ ( .D(n1941), .CLK(clk), .Q(fifo_array[290])
         );
  DFFPOSX1 fifo_array_reg_6__37_ ( .D(n1940), .CLK(clk), .Q(fifo_array[289])
         );
  DFFPOSX1 fifo_array_reg_6__36_ ( .D(n1939), .CLK(clk), .Q(fifo_array[288])
         );
  DFFPOSX1 fifo_array_reg_6__35_ ( .D(n1938), .CLK(clk), .Q(fifo_array[287])
         );
  DFFPOSX1 fifo_array_reg_6__34_ ( .D(n1937), .CLK(clk), .Q(fifo_array[286])
         );
  DFFPOSX1 fifo_array_reg_6__33_ ( .D(n1936), .CLK(clk), .Q(fifo_array[285])
         );
  DFFPOSX1 fifo_array_reg_6__32_ ( .D(n1935), .CLK(clk), .Q(fifo_array[284])
         );
  DFFPOSX1 fifo_array_reg_6__31_ ( .D(n1934), .CLK(clk), .Q(fifo_array[283])
         );
  DFFPOSX1 fifo_array_reg_6__30_ ( .D(n1933), .CLK(clk), .Q(fifo_array[282])
         );
  DFFPOSX1 fifo_array_reg_6__29_ ( .D(n1932), .CLK(clk), .Q(fifo_array[281])
         );
  DFFPOSX1 fifo_array_reg_6__28_ ( .D(n1931), .CLK(clk), .Q(fifo_array[280])
         );
  DFFPOSX1 fifo_array_reg_6__27_ ( .D(n1930), .CLK(clk), .Q(fifo_array[279])
         );
  DFFPOSX1 fifo_array_reg_6__26_ ( .D(n1929), .CLK(clk), .Q(fifo_array[278])
         );
  DFFPOSX1 fifo_array_reg_6__25_ ( .D(n1928), .CLK(clk), .Q(fifo_array[277])
         );
  DFFPOSX1 fifo_array_reg_6__24_ ( .D(n1927), .CLK(clk), .Q(fifo_array[276])
         );
  DFFPOSX1 fifo_array_reg_6__23_ ( .D(n1926), .CLK(clk), .Q(fifo_array[275])
         );
  DFFPOSX1 fifo_array_reg_6__22_ ( .D(n1925), .CLK(clk), .Q(fifo_array[274])
         );
  DFFPOSX1 fifo_array_reg_6__21_ ( .D(n1924), .CLK(clk), .Q(fifo_array[273])
         );
  DFFPOSX1 fifo_array_reg_6__20_ ( .D(n1923), .CLK(clk), .Q(fifo_array[272])
         );
  DFFPOSX1 fifo_array_reg_6__19_ ( .D(n1922), .CLK(clk), .Q(fifo_array[271])
         );
  DFFPOSX1 fifo_array_reg_6__18_ ( .D(n1921), .CLK(clk), .Q(fifo_array[270])
         );
  DFFPOSX1 fifo_array_reg_6__17_ ( .D(n1920), .CLK(clk), .Q(fifo_array[269])
         );
  DFFPOSX1 fifo_array_reg_6__16_ ( .D(n1919), .CLK(clk), .Q(fifo_array[268])
         );
  DFFPOSX1 fifo_array_reg_6__15_ ( .D(n1918), .CLK(clk), .Q(fifo_array[267])
         );
  DFFPOSX1 fifo_array_reg_6__14_ ( .D(n1917), .CLK(clk), .Q(fifo_array[266])
         );
  DFFPOSX1 fifo_array_reg_6__13_ ( .D(n1916), .CLK(clk), .Q(fifo_array[265])
         );
  DFFPOSX1 fifo_array_reg_6__12_ ( .D(n1915), .CLK(clk), .Q(fifo_array[264])
         );
  DFFPOSX1 fifo_array_reg_6__11_ ( .D(n1914), .CLK(clk), .Q(fifo_array[263])
         );
  DFFPOSX1 fifo_array_reg_6__10_ ( .D(n1913), .CLK(clk), .Q(fifo_array[262])
         );
  DFFPOSX1 fifo_array_reg_6__9_ ( .D(n1912), .CLK(clk), .Q(fifo_array[261]) );
  DFFPOSX1 fifo_array_reg_6__8_ ( .D(n1911), .CLK(clk), .Q(fifo_array[260]) );
  DFFPOSX1 fifo_array_reg_6__7_ ( .D(n1910), .CLK(clk), .Q(fifo_array[259]) );
  DFFPOSX1 fifo_array_reg_6__6_ ( .D(n1909), .CLK(clk), .Q(fifo_array[258]) );
  DFFPOSX1 fifo_array_reg_6__5_ ( .D(n1908), .CLK(clk), .Q(fifo_array[257]) );
  DFFPOSX1 fifo_array_reg_6__4_ ( .D(n1907), .CLK(clk), .Q(fifo_array[256]) );
  DFFPOSX1 fifo_array_reg_6__3_ ( .D(n1906), .CLK(clk), .Q(fifo_array[255]) );
  DFFPOSX1 fifo_array_reg_6__2_ ( .D(n1905), .CLK(clk), .Q(fifo_array[254]) );
  DFFPOSX1 fifo_array_reg_6__1_ ( .D(n1904), .CLK(clk), .Q(fifo_array[253]) );
  DFFPOSX1 fifo_array_reg_6__0_ ( .D(n1903), .CLK(clk), .Q(fifo_array[252]) );
  DFFPOSX1 fifo_array_reg_5__41_ ( .D(n1902), .CLK(clk), .Q(fifo_array[251])
         );
  DFFPOSX1 fifo_array_reg_5__40_ ( .D(n1901), .CLK(clk), .Q(fifo_array[250])
         );
  DFFPOSX1 fifo_array_reg_5__39_ ( .D(n1900), .CLK(clk), .Q(fifo_array[249])
         );
  DFFPOSX1 fifo_array_reg_5__38_ ( .D(n1899), .CLK(clk), .Q(fifo_array[248])
         );
  DFFPOSX1 fifo_array_reg_5__37_ ( .D(n1898), .CLK(clk), .Q(fifo_array[247])
         );
  DFFPOSX1 fifo_array_reg_5__36_ ( .D(n1897), .CLK(clk), .Q(fifo_array[246])
         );
  DFFPOSX1 fifo_array_reg_5__35_ ( .D(n1896), .CLK(clk), .Q(fifo_array[245])
         );
  DFFPOSX1 fifo_array_reg_5__34_ ( .D(n1895), .CLK(clk), .Q(fifo_array[244])
         );
  DFFPOSX1 fifo_array_reg_5__33_ ( .D(n1894), .CLK(clk), .Q(fifo_array[243])
         );
  DFFPOSX1 fifo_array_reg_5__32_ ( .D(n1893), .CLK(clk), .Q(fifo_array[242])
         );
  DFFPOSX1 fifo_array_reg_5__31_ ( .D(n1892), .CLK(clk), .Q(fifo_array[241])
         );
  DFFPOSX1 fifo_array_reg_5__30_ ( .D(n1891), .CLK(clk), .Q(fifo_array[240])
         );
  DFFPOSX1 fifo_array_reg_5__29_ ( .D(n1890), .CLK(clk), .Q(fifo_array[239])
         );
  DFFPOSX1 fifo_array_reg_5__28_ ( .D(n1889), .CLK(clk), .Q(fifo_array[238])
         );
  DFFPOSX1 fifo_array_reg_5__27_ ( .D(n1888), .CLK(clk), .Q(fifo_array[237])
         );
  DFFPOSX1 fifo_array_reg_5__26_ ( .D(n1887), .CLK(clk), .Q(fifo_array[236])
         );
  DFFPOSX1 fifo_array_reg_5__25_ ( .D(n1886), .CLK(clk), .Q(fifo_array[235])
         );
  DFFPOSX1 fifo_array_reg_5__24_ ( .D(n1885), .CLK(clk), .Q(fifo_array[234])
         );
  DFFPOSX1 fifo_array_reg_5__23_ ( .D(n1884), .CLK(clk), .Q(fifo_array[233])
         );
  DFFPOSX1 fifo_array_reg_5__22_ ( .D(n1883), .CLK(clk), .Q(fifo_array[232])
         );
  DFFPOSX1 fifo_array_reg_5__21_ ( .D(n1882), .CLK(clk), .Q(fifo_array[231])
         );
  DFFPOSX1 fifo_array_reg_5__20_ ( .D(n1881), .CLK(clk), .Q(fifo_array[230])
         );
  DFFPOSX1 fifo_array_reg_5__19_ ( .D(n1880), .CLK(clk), .Q(fifo_array[229])
         );
  DFFPOSX1 fifo_array_reg_5__18_ ( .D(n1879), .CLK(clk), .Q(fifo_array[228])
         );
  DFFPOSX1 fifo_array_reg_5__17_ ( .D(n1878), .CLK(clk), .Q(fifo_array[227])
         );
  DFFPOSX1 fifo_array_reg_5__16_ ( .D(n1877), .CLK(clk), .Q(fifo_array[226])
         );
  DFFPOSX1 fifo_array_reg_5__15_ ( .D(n1876), .CLK(clk), .Q(fifo_array[225])
         );
  DFFPOSX1 fifo_array_reg_5__14_ ( .D(n1875), .CLK(clk), .Q(fifo_array[224])
         );
  DFFPOSX1 fifo_array_reg_5__13_ ( .D(n1874), .CLK(clk), .Q(fifo_array[223])
         );
  DFFPOSX1 fifo_array_reg_5__12_ ( .D(n1873), .CLK(clk), .Q(fifo_array[222])
         );
  DFFPOSX1 fifo_array_reg_5__11_ ( .D(n1872), .CLK(clk), .Q(fifo_array[221])
         );
  DFFPOSX1 fifo_array_reg_5__10_ ( .D(n1871), .CLK(clk), .Q(fifo_array[220])
         );
  DFFPOSX1 fifo_array_reg_5__9_ ( .D(n1870), .CLK(clk), .Q(fifo_array[219]) );
  DFFPOSX1 fifo_array_reg_5__8_ ( .D(n1869), .CLK(clk), .Q(fifo_array[218]) );
  DFFPOSX1 fifo_array_reg_5__7_ ( .D(n1868), .CLK(clk), .Q(fifo_array[217]) );
  DFFPOSX1 fifo_array_reg_5__6_ ( .D(n1867), .CLK(clk), .Q(fifo_array[216]) );
  DFFPOSX1 fifo_array_reg_5__5_ ( .D(n1866), .CLK(clk), .Q(fifo_array[215]) );
  DFFPOSX1 fifo_array_reg_5__4_ ( .D(n1865), .CLK(clk), .Q(fifo_array[214]) );
  DFFPOSX1 fifo_array_reg_5__3_ ( .D(n1864), .CLK(clk), .Q(fifo_array[213]) );
  DFFPOSX1 fifo_array_reg_5__2_ ( .D(n1863), .CLK(clk), .Q(fifo_array[212]) );
  DFFPOSX1 fifo_array_reg_5__1_ ( .D(n1862), .CLK(clk), .Q(fifo_array[211]) );
  DFFPOSX1 fifo_array_reg_5__0_ ( .D(n1861), .CLK(clk), .Q(fifo_array[210]) );
  DFFPOSX1 fifo_array_reg_4__41_ ( .D(n1860), .CLK(clk), .Q(fifo_array[209])
         );
  DFFPOSX1 fifo_array_reg_4__40_ ( .D(n1859), .CLK(clk), .Q(fifo_array[208])
         );
  DFFPOSX1 fifo_array_reg_4__39_ ( .D(n1858), .CLK(clk), .Q(fifo_array[207])
         );
  DFFPOSX1 fifo_array_reg_4__38_ ( .D(n1857), .CLK(clk), .Q(fifo_array[206])
         );
  DFFPOSX1 fifo_array_reg_4__37_ ( .D(n1856), .CLK(clk), .Q(fifo_array[205])
         );
  DFFPOSX1 fifo_array_reg_4__36_ ( .D(n1855), .CLK(clk), .Q(fifo_array[204])
         );
  DFFPOSX1 fifo_array_reg_4__35_ ( .D(n1854), .CLK(clk), .Q(fifo_array[203])
         );
  DFFPOSX1 fifo_array_reg_4__34_ ( .D(n1853), .CLK(clk), .Q(fifo_array[202])
         );
  DFFPOSX1 fifo_array_reg_4__33_ ( .D(n1852), .CLK(clk), .Q(fifo_array[201])
         );
  DFFPOSX1 fifo_array_reg_4__32_ ( .D(n1851), .CLK(clk), .Q(fifo_array[200])
         );
  DFFPOSX1 fifo_array_reg_4__31_ ( .D(n1850), .CLK(clk), .Q(fifo_array[199])
         );
  DFFPOSX1 fifo_array_reg_4__30_ ( .D(n1849), .CLK(clk), .Q(fifo_array[198])
         );
  DFFPOSX1 fifo_array_reg_4__29_ ( .D(n1848), .CLK(clk), .Q(fifo_array[197])
         );
  DFFPOSX1 fifo_array_reg_4__28_ ( .D(n1847), .CLK(clk), .Q(fifo_array[196])
         );
  DFFPOSX1 fifo_array_reg_4__27_ ( .D(n1846), .CLK(clk), .Q(fifo_array[195])
         );
  DFFPOSX1 fifo_array_reg_4__26_ ( .D(n1845), .CLK(clk), .Q(fifo_array[194])
         );
  DFFPOSX1 fifo_array_reg_4__25_ ( .D(n1844), .CLK(clk), .Q(fifo_array[193])
         );
  DFFPOSX1 fifo_array_reg_4__24_ ( .D(n1843), .CLK(clk), .Q(fifo_array[192])
         );
  DFFPOSX1 fifo_array_reg_4__23_ ( .D(n1842), .CLK(clk), .Q(fifo_array[191])
         );
  DFFPOSX1 fifo_array_reg_4__22_ ( .D(n1841), .CLK(clk), .Q(fifo_array[190])
         );
  DFFPOSX1 fifo_array_reg_4__21_ ( .D(n1840), .CLK(clk), .Q(fifo_array[189])
         );
  DFFPOSX1 fifo_array_reg_4__20_ ( .D(n1839), .CLK(clk), .Q(fifo_array[188])
         );
  DFFPOSX1 fifo_array_reg_4__19_ ( .D(n1838), .CLK(clk), .Q(fifo_array[187])
         );
  DFFPOSX1 fifo_array_reg_4__18_ ( .D(n1837), .CLK(clk), .Q(fifo_array[186])
         );
  DFFPOSX1 fifo_array_reg_4__17_ ( .D(n1836), .CLK(clk), .Q(fifo_array[185])
         );
  DFFPOSX1 fifo_array_reg_4__16_ ( .D(n1835), .CLK(clk), .Q(fifo_array[184])
         );
  DFFPOSX1 fifo_array_reg_4__15_ ( .D(n1834), .CLK(clk), .Q(fifo_array[183])
         );
  DFFPOSX1 fifo_array_reg_4__14_ ( .D(n1833), .CLK(clk), .Q(fifo_array[182])
         );
  DFFPOSX1 fifo_array_reg_4__13_ ( .D(n1832), .CLK(clk), .Q(fifo_array[181])
         );
  DFFPOSX1 fifo_array_reg_4__12_ ( .D(n1831), .CLK(clk), .Q(fifo_array[180])
         );
  DFFPOSX1 fifo_array_reg_4__11_ ( .D(n1830), .CLK(clk), .Q(fifo_array[179])
         );
  DFFPOSX1 fifo_array_reg_4__10_ ( .D(n1829), .CLK(clk), .Q(fifo_array[178])
         );
  DFFPOSX1 fifo_array_reg_4__9_ ( .D(n1828), .CLK(clk), .Q(fifo_array[177]) );
  DFFPOSX1 fifo_array_reg_4__8_ ( .D(n1827), .CLK(clk), .Q(fifo_array[176]) );
  DFFPOSX1 fifo_array_reg_4__7_ ( .D(n1826), .CLK(clk), .Q(fifo_array[175]) );
  DFFPOSX1 fifo_array_reg_4__6_ ( .D(n1825), .CLK(clk), .Q(fifo_array[174]) );
  DFFPOSX1 fifo_array_reg_4__5_ ( .D(n1824), .CLK(clk), .Q(fifo_array[173]) );
  DFFPOSX1 fifo_array_reg_4__4_ ( .D(n1823), .CLK(clk), .Q(fifo_array[172]) );
  DFFPOSX1 fifo_array_reg_4__3_ ( .D(n1822), .CLK(clk), .Q(fifo_array[171]) );
  DFFPOSX1 fifo_array_reg_4__2_ ( .D(n1821), .CLK(clk), .Q(fifo_array[170]) );
  DFFPOSX1 fifo_array_reg_4__1_ ( .D(n1820), .CLK(clk), .Q(fifo_array[169]) );
  DFFPOSX1 fifo_array_reg_4__0_ ( .D(n1819), .CLK(clk), .Q(fifo_array[168]) );
  DFFPOSX1 fifo_array_reg_3__41_ ( .D(n1818), .CLK(clk), .Q(fifo_array[167])
         );
  DFFPOSX1 fifo_array_reg_3__40_ ( .D(n1817), .CLK(clk), .Q(fifo_array[166])
         );
  DFFPOSX1 fifo_array_reg_3__39_ ( .D(n1816), .CLK(clk), .Q(fifo_array[165])
         );
  DFFPOSX1 fifo_array_reg_3__38_ ( .D(n1815), .CLK(clk), .Q(fifo_array[164])
         );
  DFFPOSX1 fifo_array_reg_3__37_ ( .D(n1814), .CLK(clk), .Q(fifo_array[163])
         );
  DFFPOSX1 fifo_array_reg_3__36_ ( .D(n1813), .CLK(clk), .Q(fifo_array[162])
         );
  DFFPOSX1 fifo_array_reg_3__35_ ( .D(n1812), .CLK(clk), .Q(fifo_array[161])
         );
  DFFPOSX1 fifo_array_reg_3__34_ ( .D(n1811), .CLK(clk), .Q(fifo_array[160])
         );
  DFFPOSX1 fifo_array_reg_3__33_ ( .D(n1810), .CLK(clk), .Q(fifo_array[159])
         );
  DFFPOSX1 fifo_array_reg_3__32_ ( .D(n1809), .CLK(clk), .Q(fifo_array[158])
         );
  DFFPOSX1 fifo_array_reg_3__31_ ( .D(n1808), .CLK(clk), .Q(fifo_array[157])
         );
  DFFPOSX1 fifo_array_reg_3__30_ ( .D(n1807), .CLK(clk), .Q(fifo_array[156])
         );
  DFFPOSX1 fifo_array_reg_3__29_ ( .D(n1806), .CLK(clk), .Q(fifo_array[155])
         );
  DFFPOSX1 fifo_array_reg_3__28_ ( .D(n1805), .CLK(clk), .Q(fifo_array[154])
         );
  DFFPOSX1 fifo_array_reg_3__27_ ( .D(n1804), .CLK(clk), .Q(fifo_array[153])
         );
  DFFPOSX1 fifo_array_reg_3__26_ ( .D(n1803), .CLK(clk), .Q(fifo_array[152])
         );
  DFFPOSX1 fifo_array_reg_3__25_ ( .D(n1802), .CLK(clk), .Q(fifo_array[151])
         );
  DFFPOSX1 fifo_array_reg_3__24_ ( .D(n1801), .CLK(clk), .Q(fifo_array[150])
         );
  DFFPOSX1 fifo_array_reg_3__23_ ( .D(n1800), .CLK(clk), .Q(fifo_array[149])
         );
  DFFPOSX1 fifo_array_reg_3__22_ ( .D(n1799), .CLK(clk), .Q(fifo_array[148])
         );
  DFFPOSX1 fifo_array_reg_3__21_ ( .D(n1798), .CLK(clk), .Q(fifo_array[147])
         );
  DFFPOSX1 fifo_array_reg_3__20_ ( .D(n1797), .CLK(clk), .Q(fifo_array[146])
         );
  DFFPOSX1 fifo_array_reg_3__19_ ( .D(n1796), .CLK(clk), .Q(fifo_array[145])
         );
  DFFPOSX1 fifo_array_reg_3__18_ ( .D(n1795), .CLK(clk), .Q(fifo_array[144])
         );
  DFFPOSX1 fifo_array_reg_3__17_ ( .D(n1794), .CLK(clk), .Q(fifo_array[143])
         );
  DFFPOSX1 fifo_array_reg_3__16_ ( .D(n1793), .CLK(clk), .Q(fifo_array[142])
         );
  DFFPOSX1 fifo_array_reg_3__15_ ( .D(n1792), .CLK(clk), .Q(fifo_array[141])
         );
  DFFPOSX1 fifo_array_reg_3__14_ ( .D(n1791), .CLK(clk), .Q(fifo_array[140])
         );
  DFFPOSX1 fifo_array_reg_3__13_ ( .D(n1790), .CLK(clk), .Q(fifo_array[139])
         );
  DFFPOSX1 fifo_array_reg_3__12_ ( .D(n1789), .CLK(clk), .Q(fifo_array[138])
         );
  DFFPOSX1 fifo_array_reg_3__11_ ( .D(n1788), .CLK(clk), .Q(fifo_array[137])
         );
  DFFPOSX1 fifo_array_reg_3__10_ ( .D(n1787), .CLK(clk), .Q(fifo_array[136])
         );
  DFFPOSX1 fifo_array_reg_3__9_ ( .D(n1786), .CLK(clk), .Q(fifo_array[135]) );
  DFFPOSX1 fifo_array_reg_3__8_ ( .D(n1785), .CLK(clk), .Q(fifo_array[134]) );
  DFFPOSX1 fifo_array_reg_3__7_ ( .D(n1784), .CLK(clk), .Q(fifo_array[133]) );
  DFFPOSX1 fifo_array_reg_3__6_ ( .D(n1783), .CLK(clk), .Q(fifo_array[132]) );
  DFFPOSX1 fifo_array_reg_3__5_ ( .D(n1782), .CLK(clk), .Q(fifo_array[131]) );
  DFFPOSX1 fifo_array_reg_3__4_ ( .D(n1781), .CLK(clk), .Q(fifo_array[130]) );
  DFFPOSX1 fifo_array_reg_3__3_ ( .D(n1780), .CLK(clk), .Q(fifo_array[129]) );
  DFFPOSX1 fifo_array_reg_3__2_ ( .D(n1779), .CLK(clk), .Q(fifo_array[128]) );
  DFFPOSX1 fifo_array_reg_3__1_ ( .D(n1778), .CLK(clk), .Q(fifo_array[127]) );
  DFFPOSX1 fifo_array_reg_3__0_ ( .D(n1777), .CLK(clk), .Q(fifo_array[126]) );
  DFFPOSX1 fifo_array_reg_2__41_ ( .D(n1776), .CLK(clk), .Q(fifo_array[125])
         );
  DFFPOSX1 fifo_array_reg_2__40_ ( .D(n1775), .CLK(clk), .Q(fifo_array[124])
         );
  DFFPOSX1 fifo_array_reg_2__39_ ( .D(n1774), .CLK(clk), .Q(fifo_array[123])
         );
  DFFPOSX1 fifo_array_reg_2__38_ ( .D(n1773), .CLK(clk), .Q(fifo_array[122])
         );
  DFFPOSX1 fifo_array_reg_2__37_ ( .D(n1772), .CLK(clk), .Q(fifo_array[121])
         );
  DFFPOSX1 fifo_array_reg_2__36_ ( .D(n1771), .CLK(clk), .Q(fifo_array[120])
         );
  DFFPOSX1 fifo_array_reg_2__35_ ( .D(n1770), .CLK(clk), .Q(fifo_array[119])
         );
  DFFPOSX1 fifo_array_reg_2__34_ ( .D(n1769), .CLK(clk), .Q(fifo_array[118])
         );
  DFFPOSX1 fifo_array_reg_2__33_ ( .D(n1768), .CLK(clk), .Q(fifo_array[117])
         );
  DFFPOSX1 fifo_array_reg_2__32_ ( .D(n1767), .CLK(clk), .Q(fifo_array[116])
         );
  DFFPOSX1 fifo_array_reg_2__31_ ( .D(n1766), .CLK(clk), .Q(fifo_array[115])
         );
  DFFPOSX1 fifo_array_reg_2__30_ ( .D(n1765), .CLK(clk), .Q(fifo_array[114])
         );
  DFFPOSX1 fifo_array_reg_2__29_ ( .D(n1764), .CLK(clk), .Q(fifo_array[113])
         );
  DFFPOSX1 fifo_array_reg_2__28_ ( .D(n1763), .CLK(clk), .Q(fifo_array[112])
         );
  DFFPOSX1 fifo_array_reg_2__27_ ( .D(n1762), .CLK(clk), .Q(fifo_array[111])
         );
  DFFPOSX1 fifo_array_reg_2__26_ ( .D(n1761), .CLK(clk), .Q(fifo_array[110])
         );
  DFFPOSX1 fifo_array_reg_2__25_ ( .D(n1760), .CLK(clk), .Q(fifo_array[109])
         );
  DFFPOSX1 fifo_array_reg_2__24_ ( .D(n1759), .CLK(clk), .Q(fifo_array[108])
         );
  DFFPOSX1 fifo_array_reg_2__23_ ( .D(n1758), .CLK(clk), .Q(fifo_array[107])
         );
  DFFPOSX1 fifo_array_reg_2__22_ ( .D(n1757), .CLK(clk), .Q(fifo_array[106])
         );
  DFFPOSX1 fifo_array_reg_2__21_ ( .D(n1756), .CLK(clk), .Q(fifo_array[105])
         );
  DFFPOSX1 fifo_array_reg_2__20_ ( .D(n1755), .CLK(clk), .Q(fifo_array[104])
         );
  DFFPOSX1 fifo_array_reg_2__19_ ( .D(n1754), .CLK(clk), .Q(fifo_array[103])
         );
  DFFPOSX1 fifo_array_reg_2__18_ ( .D(n1753), .CLK(clk), .Q(fifo_array[102])
         );
  DFFPOSX1 fifo_array_reg_2__17_ ( .D(n1752), .CLK(clk), .Q(fifo_array[101])
         );
  DFFPOSX1 fifo_array_reg_2__16_ ( .D(n1751), .CLK(clk), .Q(fifo_array[100])
         );
  DFFPOSX1 fifo_array_reg_2__15_ ( .D(n1750), .CLK(clk), .Q(fifo_array[99]) );
  DFFPOSX1 fifo_array_reg_2__14_ ( .D(n1749), .CLK(clk), .Q(fifo_array[98]) );
  DFFPOSX1 fifo_array_reg_2__13_ ( .D(n1748), .CLK(clk), .Q(fifo_array[97]) );
  DFFPOSX1 fifo_array_reg_2__12_ ( .D(n1747), .CLK(clk), .Q(fifo_array[96]) );
  DFFPOSX1 fifo_array_reg_2__11_ ( .D(n1746), .CLK(clk), .Q(fifo_array[95]) );
  DFFPOSX1 fifo_array_reg_2__10_ ( .D(n1745), .CLK(clk), .Q(fifo_array[94]) );
  DFFPOSX1 fifo_array_reg_2__9_ ( .D(n1744), .CLK(clk), .Q(fifo_array[93]) );
  DFFPOSX1 fifo_array_reg_2__8_ ( .D(n1743), .CLK(clk), .Q(fifo_array[92]) );
  DFFPOSX1 fifo_array_reg_2__7_ ( .D(n1742), .CLK(clk), .Q(fifo_array[91]) );
  DFFPOSX1 fifo_array_reg_2__6_ ( .D(n1741), .CLK(clk), .Q(fifo_array[90]) );
  DFFPOSX1 fifo_array_reg_2__5_ ( .D(n1740), .CLK(clk), .Q(fifo_array[89]) );
  DFFPOSX1 fifo_array_reg_2__4_ ( .D(n1739), .CLK(clk), .Q(fifo_array[88]) );
  DFFPOSX1 fifo_array_reg_2__3_ ( .D(n1738), .CLK(clk), .Q(fifo_array[87]) );
  DFFPOSX1 fifo_array_reg_2__2_ ( .D(n1737), .CLK(clk), .Q(fifo_array[86]) );
  DFFPOSX1 fifo_array_reg_2__1_ ( .D(n1736), .CLK(clk), .Q(fifo_array[85]) );
  DFFPOSX1 fifo_array_reg_2__0_ ( .D(n1735), .CLK(clk), .Q(fifo_array[84]) );
  DFFPOSX1 fifo_array_reg_1__41_ ( .D(n1734), .CLK(clk), .Q(fifo_array[83]) );
  DFFPOSX1 fifo_array_reg_1__40_ ( .D(n1733), .CLK(clk), .Q(fifo_array[82]) );
  DFFPOSX1 fifo_array_reg_1__39_ ( .D(n1732), .CLK(clk), .Q(fifo_array[81]) );
  DFFPOSX1 fifo_array_reg_1__38_ ( .D(n1731), .CLK(clk), .Q(fifo_array[80]) );
  DFFPOSX1 fifo_array_reg_1__37_ ( .D(n1730), .CLK(clk), .Q(fifo_array[79]) );
  DFFPOSX1 fifo_array_reg_1__36_ ( .D(n1729), .CLK(clk), .Q(fifo_array[78]) );
  DFFPOSX1 fifo_array_reg_1__35_ ( .D(n1728), .CLK(clk), .Q(fifo_array[77]) );
  DFFPOSX1 fifo_array_reg_1__34_ ( .D(n1727), .CLK(clk), .Q(fifo_array[76]) );
  DFFPOSX1 fifo_array_reg_1__33_ ( .D(n1726), .CLK(clk), .Q(fifo_array[75]) );
  DFFPOSX1 fifo_array_reg_1__32_ ( .D(n1725), .CLK(clk), .Q(fifo_array[74]) );
  DFFPOSX1 fifo_array_reg_1__31_ ( .D(n1724), .CLK(clk), .Q(fifo_array[73]) );
  DFFPOSX1 fifo_array_reg_1__30_ ( .D(n1723), .CLK(clk), .Q(fifo_array[72]) );
  DFFPOSX1 fifo_array_reg_1__29_ ( .D(n1722), .CLK(clk), .Q(fifo_array[71]) );
  DFFPOSX1 fifo_array_reg_1__28_ ( .D(n1721), .CLK(clk), .Q(fifo_array[70]) );
  DFFPOSX1 fifo_array_reg_1__27_ ( .D(n1720), .CLK(clk), .Q(fifo_array[69]) );
  DFFPOSX1 fifo_array_reg_1__26_ ( .D(n1719), .CLK(clk), .Q(fifo_array[68]) );
  DFFPOSX1 fifo_array_reg_1__25_ ( .D(n1718), .CLK(clk), .Q(fifo_array[67]) );
  DFFPOSX1 fifo_array_reg_1__24_ ( .D(n1717), .CLK(clk), .Q(fifo_array[66]) );
  DFFPOSX1 fifo_array_reg_1__23_ ( .D(n1716), .CLK(clk), .Q(fifo_array[65]) );
  DFFPOSX1 fifo_array_reg_1__22_ ( .D(n1715), .CLK(clk), .Q(fifo_array[64]) );
  DFFPOSX1 fifo_array_reg_1__21_ ( .D(n1714), .CLK(clk), .Q(fifo_array[63]) );
  DFFPOSX1 fifo_array_reg_1__20_ ( .D(n1713), .CLK(clk), .Q(fifo_array[62]) );
  DFFPOSX1 fifo_array_reg_1__19_ ( .D(n1712), .CLK(clk), .Q(fifo_array[61]) );
  DFFPOSX1 fifo_array_reg_1__18_ ( .D(n1711), .CLK(clk), .Q(fifo_array[60]) );
  DFFPOSX1 fifo_array_reg_1__17_ ( .D(n1710), .CLK(clk), .Q(fifo_array[59]) );
  DFFPOSX1 fifo_array_reg_1__16_ ( .D(n1709), .CLK(clk), .Q(fifo_array[58]) );
  DFFPOSX1 fifo_array_reg_1__15_ ( .D(n1708), .CLK(clk), .Q(fifo_array[57]) );
  DFFPOSX1 fifo_array_reg_1__14_ ( .D(n1707), .CLK(clk), .Q(fifo_array[56]) );
  DFFPOSX1 fifo_array_reg_1__13_ ( .D(n1706), .CLK(clk), .Q(fifo_array[55]) );
  DFFPOSX1 fifo_array_reg_1__12_ ( .D(n1705), .CLK(clk), .Q(fifo_array[54]) );
  DFFPOSX1 fifo_array_reg_1__11_ ( .D(n1704), .CLK(clk), .Q(fifo_array[53]) );
  DFFPOSX1 fifo_array_reg_1__10_ ( .D(n1703), .CLK(clk), .Q(fifo_array[52]) );
  DFFPOSX1 fifo_array_reg_1__9_ ( .D(n1702), .CLK(clk), .Q(fifo_array[51]) );
  DFFPOSX1 fifo_array_reg_1__8_ ( .D(n1701), .CLK(clk), .Q(fifo_array[50]) );
  DFFPOSX1 fifo_array_reg_1__7_ ( .D(n1700), .CLK(clk), .Q(fifo_array[49]) );
  DFFPOSX1 fifo_array_reg_1__6_ ( .D(n1699), .CLK(clk), .Q(fifo_array[48]) );
  DFFPOSX1 fifo_array_reg_1__5_ ( .D(n1698), .CLK(clk), .Q(fifo_array[47]) );
  DFFPOSX1 fifo_array_reg_1__4_ ( .D(n1697), .CLK(clk), .Q(fifo_array[46]) );
  DFFPOSX1 fifo_array_reg_1__3_ ( .D(n1696), .CLK(clk), .Q(fifo_array[45]) );
  DFFPOSX1 fifo_array_reg_1__2_ ( .D(n1695), .CLK(clk), .Q(fifo_array[44]) );
  DFFPOSX1 fifo_array_reg_1__1_ ( .D(n1694), .CLK(clk), .Q(fifo_array[43]) );
  DFFPOSX1 fifo_array_reg_1__0_ ( .D(n1693), .CLK(clk), .Q(fifo_array[42]) );
  DFFPOSX1 fifo_array_reg_0__41_ ( .D(n1692), .CLK(clk), .Q(fifo_array[41]) );
  DFFPOSX1 fifo_array_reg_0__40_ ( .D(n1691), .CLK(clk), .Q(fifo_array[40]) );
  DFFPOSX1 fifo_array_reg_0__39_ ( .D(n1690), .CLK(clk), .Q(fifo_array[39]) );
  DFFPOSX1 fifo_array_reg_0__38_ ( .D(n1689), .CLK(clk), .Q(fifo_array[38]) );
  DFFPOSX1 fifo_array_reg_0__37_ ( .D(n1688), .CLK(clk), .Q(fifo_array[37]) );
  DFFPOSX1 fifo_array_reg_0__36_ ( .D(n1687), .CLK(clk), .Q(fifo_array[36]) );
  DFFPOSX1 fifo_array_reg_0__35_ ( .D(n1686), .CLK(clk), .Q(fifo_array[35]) );
  DFFPOSX1 fifo_array_reg_0__34_ ( .D(n1685), .CLK(clk), .Q(fifo_array[34]) );
  DFFPOSX1 fifo_array_reg_0__33_ ( .D(n1684), .CLK(clk), .Q(fifo_array[33]) );
  DFFPOSX1 fifo_array_reg_0__32_ ( .D(n1683), .CLK(clk), .Q(fifo_array[32]) );
  DFFPOSX1 fifo_array_reg_0__31_ ( .D(n1682), .CLK(clk), .Q(fifo_array[31]) );
  DFFPOSX1 fifo_array_reg_0__30_ ( .D(n1681), .CLK(clk), .Q(fifo_array[30]) );
  DFFPOSX1 fifo_array_reg_0__29_ ( .D(n1680), .CLK(clk), .Q(fifo_array[29]) );
  DFFPOSX1 fifo_array_reg_0__28_ ( .D(n1679), .CLK(clk), .Q(fifo_array[28]) );
  DFFPOSX1 fifo_array_reg_0__27_ ( .D(n1678), .CLK(clk), .Q(fifo_array[27]) );
  DFFPOSX1 fifo_array_reg_0__26_ ( .D(n1677), .CLK(clk), .Q(fifo_array[26]) );
  DFFPOSX1 fifo_array_reg_0__25_ ( .D(n1676), .CLK(clk), .Q(fifo_array[25]) );
  DFFPOSX1 fifo_array_reg_0__24_ ( .D(n1675), .CLK(clk), .Q(fifo_array[24]) );
  DFFPOSX1 fifo_array_reg_0__23_ ( .D(n1674), .CLK(clk), .Q(fifo_array[23]) );
  DFFPOSX1 fifo_array_reg_0__22_ ( .D(n1673), .CLK(clk), .Q(fifo_array[22]) );
  DFFPOSX1 fifo_array_reg_0__21_ ( .D(n1672), .CLK(clk), .Q(fifo_array[21]) );
  DFFPOSX1 fifo_array_reg_0__20_ ( .D(n1671), .CLK(clk), .Q(fifo_array[20]) );
  DFFPOSX1 fifo_array_reg_0__19_ ( .D(n1670), .CLK(clk), .Q(fifo_array[19]) );
  DFFPOSX1 fifo_array_reg_0__18_ ( .D(n1669), .CLK(clk), .Q(fifo_array[18]) );
  DFFPOSX1 fifo_array_reg_0__17_ ( .D(n1668), .CLK(clk), .Q(fifo_array[17]) );
  DFFPOSX1 fifo_array_reg_0__16_ ( .D(n1667), .CLK(clk), .Q(fifo_array[16]) );
  DFFPOSX1 fifo_array_reg_0__15_ ( .D(n1666), .CLK(clk), .Q(fifo_array[15]) );
  DFFPOSX1 fifo_array_reg_0__14_ ( .D(n1665), .CLK(clk), .Q(fifo_array[14]) );
  DFFPOSX1 fifo_array_reg_0__13_ ( .D(n1664), .CLK(clk), .Q(fifo_array[13]) );
  DFFPOSX1 fifo_array_reg_0__12_ ( .D(n1663), .CLK(clk), .Q(fifo_array[12]) );
  DFFPOSX1 fifo_array_reg_0__11_ ( .D(n1662), .CLK(clk), .Q(fifo_array[11]) );
  DFFPOSX1 fifo_array_reg_0__10_ ( .D(n1661), .CLK(clk), .Q(fifo_array[10]) );
  DFFPOSX1 fifo_array_reg_0__9_ ( .D(n1660), .CLK(clk), .Q(fifo_array[9]) );
  DFFPOSX1 fifo_array_reg_0__8_ ( .D(n1659), .CLK(clk), .Q(fifo_array[8]) );
  DFFPOSX1 fifo_array_reg_0__7_ ( .D(n1658), .CLK(clk), .Q(fifo_array[7]) );
  DFFPOSX1 fifo_array_reg_0__6_ ( .D(n1657), .CLK(clk), .Q(fifo_array[6]) );
  DFFPOSX1 fifo_array_reg_0__5_ ( .D(n1656), .CLK(clk), .Q(fifo_array[5]) );
  DFFPOSX1 fifo_array_reg_0__4_ ( .D(n1655), .CLK(clk), .Q(fifo_array[4]) );
  DFFPOSX1 fifo_array_reg_0__3_ ( .D(n1654), .CLK(clk), .Q(fifo_array[3]) );
  DFFPOSX1 fifo_array_reg_0__2_ ( .D(n1653), .CLK(clk), .Q(fifo_array[2]) );
  DFFPOSX1 fifo_array_reg_0__1_ ( .D(n1652), .CLK(clk), .Q(fifo_array[1]) );
  DFFPOSX1 fifo_array_reg_0__0_ ( .D(n1651), .CLK(clk), .Q(fifo_array[0]) );
  OAI21X1 U118 ( .A(n5839), .B(n5746), .C(n4317), .Y(n1651) );
  OAI21X1 U120 ( .A(n5838), .B(n5745), .C(n4226), .Y(n1652) );
  OAI21X1 U122 ( .A(n5838), .B(n5744), .C(n4138), .Y(n1653) );
  OAI21X1 U124 ( .A(n5838), .B(n5743), .C(n4049), .Y(n1654) );
  OAI21X1 U126 ( .A(n5838), .B(n5742), .C(n3956), .Y(n1655) );
  OAI21X1 U128 ( .A(n5838), .B(n5741), .C(n3874), .Y(n1656) );
  OAI21X1 U130 ( .A(n5838), .B(n5740), .C(n3791), .Y(n1657) );
  OAI21X1 U132 ( .A(n5838), .B(n5739), .C(n3709), .Y(n1658) );
  OAI21X1 U134 ( .A(n5838), .B(n5738), .C(n4316), .Y(n1659) );
  OAI21X1 U136 ( .A(n5838), .B(n5737), .C(n3628), .Y(n1660) );
  OAI21X1 U138 ( .A(n5838), .B(n5736), .C(n3551), .Y(n1661) );
  OAI21X1 U140 ( .A(n5838), .B(n5735), .C(n3472), .Y(n1662) );
  OAI21X1 U142 ( .A(n5838), .B(n5734), .C(n3394), .Y(n1663) );
  OAI21X1 U144 ( .A(n5838), .B(n5733), .C(n4225), .Y(n1664) );
  OAI21X1 U146 ( .A(n5838), .B(n5732), .C(n4137), .Y(n1665) );
  OAI21X1 U148 ( .A(n5839), .B(n5731), .C(n4048), .Y(n1666) );
  OAI21X1 U150 ( .A(n5838), .B(n5749), .C(n3627), .Y(n1667) );
  OAI21X1 U152 ( .A(n5839), .B(n5750), .C(n3955), .Y(n1668) );
  OAI21X1 U154 ( .A(n5838), .B(n5751), .C(n3873), .Y(n1669) );
  OAI21X1 U156 ( .A(n5839), .B(n5752), .C(n3790), .Y(n1670) );
  OAI21X1 U158 ( .A(n5839), .B(n5753), .C(n3708), .Y(n1671) );
  OAI21X1 U160 ( .A(n5838), .B(n5754), .C(n4315), .Y(n1672) );
  OAI21X1 U162 ( .A(n5838), .B(n5755), .C(n3550), .Y(n1673) );
  OAI21X1 U164 ( .A(n5838), .B(n5756), .C(n3471), .Y(n1674) );
  OAI21X1 U166 ( .A(n5838), .B(n5757), .C(n3393), .Y(n1675) );
  OAI21X1 U168 ( .A(n5839), .B(n5758), .C(n4224), .Y(n1676) );
  OAI21X1 U170 ( .A(n5838), .B(n5759), .C(n4136), .Y(n1677) );
  OAI21X1 U172 ( .A(n5839), .B(n5760), .C(n3872), .Y(n1678) );
  OAI21X1 U174 ( .A(n5838), .B(n5761), .C(n3789), .Y(n1679) );
  OAI21X1 U176 ( .A(n5839), .B(n5762), .C(n3707), .Y(n1680) );
  OAI21X1 U178 ( .A(n5838), .B(n5763), .C(n3392), .Y(n1681) );
  OAI21X1 U180 ( .A(n5839), .B(n5764), .C(n3316), .Y(n1682) );
  OAI21X1 U182 ( .A(n5838), .B(n5765), .C(n3240), .Y(n1683) );
  OAI21X1 U184 ( .A(n5838), .B(n5766), .C(n3164), .Y(n1684) );
  OAI21X1 U186 ( .A(n5839), .B(n5767), .C(n3087), .Y(n1685) );
  OAI21X1 U188 ( .A(n5839), .B(n5768), .C(n1585), .Y(n1686) );
  OAI21X1 U190 ( .A(n5839), .B(n5769), .C(n3549), .Y(n1687) );
  OAI21X1 U192 ( .A(n5839), .B(n5770), .C(n3315), .Y(n1688) );
  OAI21X1 U194 ( .A(n5839), .B(n5771), .C(n3239), .Y(n1689) );
  OAI21X1 U196 ( .A(n5838), .B(n5772), .C(n3470), .Y(n1690) );
  OAI21X1 U198 ( .A(n5838), .B(n5748), .C(n3086), .Y(n1691) );
  OAI21X1 U200 ( .A(n5838), .B(n5747), .C(n177), .Y(n1692) );
  OAI21X1 U203 ( .A(n5746), .B(n5837), .C(n4223), .Y(n1693) );
  OAI21X1 U205 ( .A(n5745), .B(n5836), .C(n4314), .Y(n1694) );
  OAI21X1 U207 ( .A(n5744), .B(n5837), .C(n4047), .Y(n1695) );
  OAI21X1 U209 ( .A(n5743), .B(n5837), .C(n4135), .Y(n1696) );
  OAI21X1 U211 ( .A(n5742), .B(n5837), .C(n3871), .Y(n1697) );
  OAI21X1 U213 ( .A(n5741), .B(n5836), .C(n3954), .Y(n1698) );
  OAI21X1 U215 ( .A(n5740), .B(n5836), .C(n3706), .Y(n1699) );
  OAI21X1 U217 ( .A(n5739), .B(n5836), .C(n3788), .Y(n1700) );
  OAI21X1 U219 ( .A(n5738), .B(n5837), .C(n4222), .Y(n1701) );
  OAI21X1 U221 ( .A(n5737), .B(n5836), .C(n3548), .Y(n1702) );
  OAI21X1 U223 ( .A(n5736), .B(n5836), .C(n3626), .Y(n1703) );
  OAI21X1 U225 ( .A(n5735), .B(n5837), .C(n3391), .Y(n1704) );
  OAI21X1 U227 ( .A(n5734), .B(n5836), .C(n3469), .Y(n1705) );
  OAI21X1 U229 ( .A(n5733), .B(n5836), .C(n4313), .Y(n1706) );
  OAI21X1 U231 ( .A(n5732), .B(n5837), .C(n4046), .Y(n1707) );
  OAI21X1 U233 ( .A(n5731), .B(n5836), .C(n4134), .Y(n1708) );
  OAI21X1 U235 ( .A(n5749), .B(n5837), .C(n3547), .Y(n1709) );
  OAI21X1 U237 ( .A(n5750), .B(n5836), .C(n3870), .Y(n1710) );
  OAI21X1 U239 ( .A(n5751), .B(n5837), .C(n3953), .Y(n1711) );
  OAI21X1 U241 ( .A(n5752), .B(n5836), .C(n3705), .Y(n1712) );
  OAI21X1 U243 ( .A(n5753), .B(n5837), .C(n3787), .Y(n1713) );
  OAI21X1 U245 ( .A(n5754), .B(n5836), .C(n4221), .Y(n1714) );
  OAI21X1 U247 ( .A(n5755), .B(n5836), .C(n3625), .Y(n1715) );
  OAI21X1 U249 ( .A(n5756), .B(n5837), .C(n3390), .Y(n1716) );
  OAI21X1 U251 ( .A(n5757), .B(n5837), .C(n3468), .Y(n1717) );
  OAI21X1 U253 ( .A(n5758), .B(n5837), .C(n4312), .Y(n1718) );
  OAI21X1 U255 ( .A(n5759), .B(n5837), .C(n4045), .Y(n1719) );
  OAI21X1 U257 ( .A(n5760), .B(n5836), .C(n3952), .Y(n1720) );
  OAI21X1 U259 ( .A(n5761), .B(n5836), .C(n3704), .Y(n1721) );
  OAI21X1 U261 ( .A(n5762), .B(n5837), .C(n3786), .Y(n1722) );
  OAI21X1 U263 ( .A(n5763), .B(n5837), .C(n3467), .Y(n1723) );
  OAI21X1 U265 ( .A(n5764), .B(n5836), .C(n3238), .Y(n1724) );
  OAI21X1 U267 ( .A(n5765), .B(n5836), .C(n3314), .Y(n1725) );
  OAI21X1 U269 ( .A(n5766), .B(n5836), .C(n3085), .Y(n1726) );
  OAI21X1 U271 ( .A(n5767), .B(n5837), .C(n3163), .Y(n1727) );
  OAI21X1 U273 ( .A(n5768), .B(n5836), .C(n176), .Y(n1728) );
  OAI21X1 U275 ( .A(n5769), .B(n5837), .C(n3624), .Y(n1729) );
  OAI21X1 U277 ( .A(n5770), .B(n5836), .C(n3237), .Y(n1730) );
  OAI21X1 U279 ( .A(n5771), .B(n5836), .C(n3313), .Y(n1731) );
  OAI21X1 U281 ( .A(n5772), .B(n5836), .C(n3389), .Y(n1732) );
  OAI21X1 U283 ( .A(n5748), .B(n5836), .C(n3162), .Y(n1733) );
  OAI21X1 U285 ( .A(n5747), .B(n5836), .C(n175), .Y(n1734) );
  OAI21X1 U288 ( .A(n5746), .B(n5835), .C(n4133), .Y(n1735) );
  OAI21X1 U290 ( .A(n5745), .B(n5834), .C(n4044), .Y(n1736) );
  OAI21X1 U292 ( .A(n5744), .B(n5835), .C(n4311), .Y(n1737) );
  OAI21X1 U294 ( .A(n5743), .B(n5835), .C(n4220), .Y(n1738) );
  OAI21X1 U296 ( .A(n5742), .B(n5835), .C(n3785), .Y(n1739) );
  OAI21X1 U298 ( .A(n5741), .B(n5834), .C(n3703), .Y(n1740) );
  OAI21X1 U300 ( .A(n5740), .B(n5834), .C(n3951), .Y(n1741) );
  OAI21X1 U302 ( .A(n5739), .B(n5834), .C(n3869), .Y(n1742) );
  OAI21X1 U304 ( .A(n5738), .B(n5835), .C(n4132), .Y(n1743) );
  OAI21X1 U306 ( .A(n5737), .B(n5834), .C(n3466), .Y(n1744) );
  OAI21X1 U308 ( .A(n5736), .B(n5834), .C(n3388), .Y(n1745) );
  OAI21X1 U310 ( .A(n5735), .B(n5835), .C(n3623), .Y(n1746) );
  OAI21X1 U312 ( .A(n5734), .B(n5834), .C(n3546), .Y(n1747) );
  OAI21X1 U314 ( .A(n5733), .B(n5834), .C(n4043), .Y(n1748) );
  OAI21X1 U316 ( .A(n5732), .B(n5835), .C(n4310), .Y(n1749) );
  OAI21X1 U318 ( .A(n5731), .B(n5834), .C(n4219), .Y(n1750) );
  OAI21X1 U320 ( .A(n5749), .B(n5835), .C(n3465), .Y(n1751) );
  OAI21X1 U322 ( .A(n5750), .B(n5834), .C(n3784), .Y(n1752) );
  OAI21X1 U324 ( .A(n5751), .B(n5835), .C(n3702), .Y(n1753) );
  OAI21X1 U326 ( .A(n5752), .B(n5834), .C(n3950), .Y(n1754) );
  OAI21X1 U328 ( .A(n5753), .B(n5835), .C(n3868), .Y(n1755) );
  OAI21X1 U330 ( .A(n5754), .B(n5834), .C(n4131), .Y(n1756) );
  OAI21X1 U332 ( .A(n5755), .B(n5834), .C(n3387), .Y(n1757) );
  OAI21X1 U334 ( .A(n5756), .B(n5835), .C(n3622), .Y(n1758) );
  OAI21X1 U336 ( .A(n5757), .B(n5835), .C(n3545), .Y(n1759) );
  OAI21X1 U338 ( .A(n5758), .B(n5835), .C(n4042), .Y(n1760) );
  OAI21X1 U340 ( .A(n5759), .B(n5835), .C(n4309), .Y(n1761) );
  OAI21X1 U342 ( .A(n5760), .B(n5834), .C(n3701), .Y(n1762) );
  OAI21X1 U344 ( .A(n5761), .B(n5834), .C(n3949), .Y(n1763) );
  OAI21X1 U346 ( .A(n5762), .B(n5835), .C(n3867), .Y(n1764) );
  OAI21X1 U348 ( .A(n5763), .B(n5835), .C(n3544), .Y(n1765) );
  OAI21X1 U350 ( .A(n5764), .B(n5834), .C(n3161), .Y(n1766) );
  OAI21X1 U352 ( .A(n5765), .B(n5834), .C(n3084), .Y(n1767) );
  OAI21X1 U354 ( .A(n5766), .B(n5834), .C(n3312), .Y(n1768) );
  OAI21X1 U356 ( .A(n5767), .B(n5835), .C(n3236), .Y(n1769) );
  OAI21X1 U358 ( .A(n5768), .B(n5834), .C(n174), .Y(n1770) );
  OAI21X1 U360 ( .A(n5769), .B(n5835), .C(n3386), .Y(n1771) );
  OAI21X1 U362 ( .A(n5770), .B(n5834), .C(n3160), .Y(n1772) );
  OAI21X1 U364 ( .A(n5771), .B(n5834), .C(n3083), .Y(n1773) );
  OAI21X1 U366 ( .A(n5772), .B(n5834), .C(n3621), .Y(n1774) );
  OAI21X1 U368 ( .A(n5748), .B(n5834), .C(n3235), .Y(n1775) );
  OAI21X1 U370 ( .A(n5747), .B(n5834), .C(n173), .Y(n1776) );
  OAI21X1 U373 ( .A(n5746), .B(n5833), .C(n4041), .Y(n1777) );
  OAI21X1 U375 ( .A(n5745), .B(n5832), .C(n4130), .Y(n1778) );
  OAI21X1 U377 ( .A(n5744), .B(n5833), .C(n4218), .Y(n1779) );
  OAI21X1 U379 ( .A(n5743), .B(n5833), .C(n4308), .Y(n1780) );
  OAI21X1 U381 ( .A(n5742), .B(n5833), .C(n3700), .Y(n1781) );
  OAI21X1 U383 ( .A(n5741), .B(n5832), .C(n3783), .Y(n1782) );
  OAI21X1 U385 ( .A(n5740), .B(n5832), .C(n3866), .Y(n1783) );
  OAI21X1 U387 ( .A(n5739), .B(n5832), .C(n3948), .Y(n1784) );
  OAI21X1 U389 ( .A(n5738), .B(n5833), .C(n4040), .Y(n1785) );
  OAI21X1 U391 ( .A(n5737), .B(n5832), .C(n3385), .Y(n1786) );
  OAI21X1 U393 ( .A(n5736), .B(n5832), .C(n3464), .Y(n1787) );
  OAI21X1 U395 ( .A(n5735), .B(n5833), .C(n3543), .Y(n1788) );
  OAI21X1 U397 ( .A(n5734), .B(n5832), .C(n3620), .Y(n1789) );
  OAI21X1 U399 ( .A(n5733), .B(n5832), .C(n4129), .Y(n1790) );
  OAI21X1 U401 ( .A(n5732), .B(n5833), .C(n4217), .Y(n1791) );
  OAI21X1 U403 ( .A(n5731), .B(n5832), .C(n4307), .Y(n1792) );
  OAI21X1 U405 ( .A(n5749), .B(n5833), .C(n3384), .Y(n1793) );
  OAI21X1 U407 ( .A(n5750), .B(n5832), .C(n3699), .Y(n1794) );
  OAI21X1 U409 ( .A(n5751), .B(n5833), .C(n3782), .Y(n1795) );
  OAI21X1 U411 ( .A(n5752), .B(n5832), .C(n3865), .Y(n1796) );
  OAI21X1 U413 ( .A(n5753), .B(n5833), .C(n3947), .Y(n1797) );
  OAI21X1 U415 ( .A(n5754), .B(n5832), .C(n4039), .Y(n1798) );
  OAI21X1 U417 ( .A(n5755), .B(n5832), .C(n3463), .Y(n1799) );
  OAI21X1 U419 ( .A(n5756), .B(n5833), .C(n3542), .Y(n1800) );
  OAI21X1 U421 ( .A(n5757), .B(n5833), .C(n3619), .Y(n1801) );
  OAI21X1 U423 ( .A(n5758), .B(n5833), .C(n4128), .Y(n1802) );
  OAI21X1 U425 ( .A(n5759), .B(n5833), .C(n4216), .Y(n1803) );
  OAI21X1 U427 ( .A(n5760), .B(n5832), .C(n3781), .Y(n1804) );
  OAI21X1 U429 ( .A(n5761), .B(n5832), .C(n3864), .Y(n1805) );
  OAI21X1 U431 ( .A(n5762), .B(n5833), .C(n3946), .Y(n1806) );
  OAI21X1 U433 ( .A(n5763), .B(n5833), .C(n3618), .Y(n1807) );
  OAI21X1 U435 ( .A(n5764), .B(n5832), .C(n3082), .Y(n1808) );
  OAI21X1 U437 ( .A(n5765), .B(n5832), .C(n3159), .Y(n1809) );
  OAI21X1 U439 ( .A(n5766), .B(n5832), .C(n3234), .Y(n1810) );
  OAI21X1 U441 ( .A(n5767), .B(n5833), .C(n3311), .Y(n1811) );
  OAI21X1 U443 ( .A(n5768), .B(n5832), .C(n172), .Y(n1812) );
  OAI21X1 U445 ( .A(n5769), .B(n5833), .C(n3462), .Y(n1813) );
  OAI21X1 U447 ( .A(n5770), .B(n5832), .C(n3081), .Y(n1814) );
  OAI21X1 U449 ( .A(n5771), .B(n5832), .C(n3158), .Y(n1815) );
  OAI21X1 U451 ( .A(n5772), .B(n5832), .C(n3541), .Y(n1816) );
  OAI21X1 U453 ( .A(n5748), .B(n5832), .C(n3310), .Y(n1817) );
  OAI21X1 U455 ( .A(n5747), .B(n5832), .C(n171), .Y(n1818) );
  OAI21X1 U458 ( .A(n5746), .B(n5831), .C(n3945), .Y(n1819) );
  OAI21X1 U460 ( .A(n5745), .B(n5830), .C(n3863), .Y(n1820) );
  OAI21X1 U462 ( .A(n5744), .B(n5831), .C(n3780), .Y(n1821) );
  OAI21X1 U464 ( .A(n5743), .B(n5831), .C(n3698), .Y(n1822) );
  OAI21X1 U466 ( .A(n5742), .B(n5831), .C(n4306), .Y(n1823) );
  OAI21X1 U468 ( .A(n5741), .B(n5830), .C(n4215), .Y(n1824) );
  OAI21X1 U470 ( .A(n5740), .B(n5830), .C(n4127), .Y(n1825) );
  OAI21X1 U472 ( .A(n5739), .B(n5830), .C(n4038), .Y(n1826) );
  OAI21X1 U474 ( .A(n5738), .B(n5831), .C(n3944), .Y(n1827) );
  OAI21X1 U476 ( .A(n5737), .B(n5830), .C(n3309), .Y(n1828) );
  OAI21X1 U478 ( .A(n5736), .B(n5830), .C(n3233), .Y(n1829) );
  OAI21X1 U480 ( .A(n5735), .B(n5831), .C(n3157), .Y(n1830) );
  OAI21X1 U482 ( .A(n5734), .B(n5830), .C(n3080), .Y(n1831) );
  OAI21X1 U484 ( .A(n5733), .B(n5830), .C(n3862), .Y(n1832) );
  OAI21X1 U486 ( .A(n5732), .B(n5831), .C(n3779), .Y(n1833) );
  OAI21X1 U488 ( .A(n5731), .B(n5830), .C(n3697), .Y(n1834) );
  OAI21X1 U490 ( .A(n5749), .B(n5831), .C(n3308), .Y(n1835) );
  OAI21X1 U492 ( .A(n5750), .B(n5830), .C(n4305), .Y(n1836) );
  OAI21X1 U494 ( .A(n5751), .B(n5831), .C(n4214), .Y(n1837) );
  OAI21X1 U496 ( .A(n5752), .B(n5830), .C(n4126), .Y(n1838) );
  OAI21X1 U498 ( .A(n5753), .B(n5831), .C(n4037), .Y(n1839) );
  OAI21X1 U500 ( .A(n5754), .B(n5830), .C(n3943), .Y(n1840) );
  OAI21X1 U502 ( .A(n5755), .B(n5830), .C(n3232), .Y(n1841) );
  OAI21X1 U504 ( .A(n5756), .B(n5831), .C(n3156), .Y(n1842) );
  OAI21X1 U506 ( .A(n5757), .B(n5831), .C(n3079), .Y(n1843) );
  OAI21X1 U508 ( .A(n5758), .B(n5831), .C(n3861), .Y(n1844) );
  OAI21X1 U510 ( .A(n5759), .B(n5831), .C(n3778), .Y(n1845) );
  OAI21X1 U512 ( .A(n5760), .B(n5830), .C(n4213), .Y(n1846) );
  OAI21X1 U514 ( .A(n5761), .B(n5830), .C(n4125), .Y(n1847) );
  OAI21X1 U516 ( .A(n5762), .B(n5831), .C(n4036), .Y(n1848) );
  OAI21X1 U518 ( .A(n5763), .B(n5831), .C(n3078), .Y(n1849) );
  OAI21X1 U520 ( .A(n5764), .B(n5830), .C(n3617), .Y(n1850) );
  OAI21X1 U522 ( .A(n5765), .B(n5830), .C(n3540), .Y(n1851) );
  OAI21X1 U524 ( .A(n5766), .B(n5830), .C(n3461), .Y(n1852) );
  OAI21X1 U526 ( .A(n5767), .B(n5831), .C(n3383), .Y(n1853) );
  OAI21X1 U528 ( .A(n5768), .B(n5830), .C(n170), .Y(n1854) );
  OAI21X1 U530 ( .A(n5769), .B(n5831), .C(n3231), .Y(n1855) );
  OAI21X1 U532 ( .A(n5770), .B(n5830), .C(n3616), .Y(n1856) );
  OAI21X1 U534 ( .A(n5771), .B(n5830), .C(n3539), .Y(n1857) );
  OAI21X1 U536 ( .A(n5772), .B(n5830), .C(n3155), .Y(n1858) );
  OAI21X1 U538 ( .A(n5748), .B(n5830), .C(n3382), .Y(n1859) );
  OAI21X1 U540 ( .A(n5747), .B(n5830), .C(n169), .Y(n1860) );
  OAI21X1 U543 ( .A(n5746), .B(n5829), .C(n3860), .Y(n1861) );
  OAI21X1 U545 ( .A(n5745), .B(n5828), .C(n3942), .Y(n1862) );
  OAI21X1 U547 ( .A(n5744), .B(n5829), .C(n3696), .Y(n1863) );
  OAI21X1 U549 ( .A(n5743), .B(n5829), .C(n3777), .Y(n1864) );
  OAI21X1 U551 ( .A(n5742), .B(n5829), .C(n4212), .Y(n1865) );
  OAI21X1 U553 ( .A(n5741), .B(n5828), .C(n4304), .Y(n1866) );
  OAI21X1 U555 ( .A(n5740), .B(n5828), .C(n4035), .Y(n1867) );
  OAI21X1 U557 ( .A(n5739), .B(n5828), .C(n4124), .Y(n1868) );
  OAI21X1 U559 ( .A(n5738), .B(n5829), .C(n3859), .Y(n1869) );
  OAI21X1 U561 ( .A(n5737), .B(n5828), .C(n3230), .Y(n1870) );
  OAI21X1 U563 ( .A(n5736), .B(n5828), .C(n3307), .Y(n1871) );
  OAI21X1 U565 ( .A(n5735), .B(n5829), .C(n3077), .Y(n1872) );
  OAI21X1 U567 ( .A(n5734), .B(n5828), .C(n3154), .Y(n1873) );
  OAI21X1 U569 ( .A(n5733), .B(n5828), .C(n3941), .Y(n1874) );
  OAI21X1 U571 ( .A(n5732), .B(n5829), .C(n3695), .Y(n1875) );
  OAI21X1 U573 ( .A(n5731), .B(n5828), .C(n3776), .Y(n1876) );
  OAI21X1 U575 ( .A(n5749), .B(n5829), .C(n3229), .Y(n1877) );
  OAI21X1 U577 ( .A(n5750), .B(n5828), .C(n4211), .Y(n1878) );
  OAI21X1 U579 ( .A(n5751), .B(n5829), .C(n4303), .Y(n1879) );
  OAI21X1 U581 ( .A(n5752), .B(n5828), .C(n4034), .Y(n1880) );
  OAI21X1 U583 ( .A(n5753), .B(n5829), .C(n4123), .Y(n1881) );
  OAI21X1 U585 ( .A(n5754), .B(n5828), .C(n3858), .Y(n1882) );
  OAI21X1 U587 ( .A(n5755), .B(n5828), .C(n3306), .Y(n1883) );
  OAI21X1 U589 ( .A(n5756), .B(n5829), .C(n3076), .Y(n1884) );
  OAI21X1 U591 ( .A(n5757), .B(n5829), .C(n3153), .Y(n1885) );
  OAI21X1 U593 ( .A(n5758), .B(n5829), .C(n3940), .Y(n1886) );
  OAI21X1 U595 ( .A(n5759), .B(n5829), .C(n3694), .Y(n1887) );
  OAI21X1 U597 ( .A(n5760), .B(n5828), .C(n4302), .Y(n1888) );
  OAI21X1 U599 ( .A(n5761), .B(n5828), .C(n4033), .Y(n1889) );
  OAI21X1 U601 ( .A(n5762), .B(n5829), .C(n4122), .Y(n1890) );
  OAI21X1 U603 ( .A(n5763), .B(n5829), .C(n3152), .Y(n1891) );
  OAI21X1 U605 ( .A(n5764), .B(n5828), .C(n3538), .Y(n1892) );
  OAI21X1 U607 ( .A(n5765), .B(n5828), .C(n3615), .Y(n1893) );
  OAI21X1 U609 ( .A(n5766), .B(n5828), .C(n3381), .Y(n1894) );
  OAI21X1 U611 ( .A(n5767), .B(n5829), .C(n3460), .Y(n1895) );
  OAI21X1 U613 ( .A(n5768), .B(n5828), .C(n168), .Y(n1896) );
  OAI21X1 U615 ( .A(n5769), .B(n5829), .C(n3305), .Y(n1897) );
  OAI21X1 U617 ( .A(n5770), .B(n5828), .C(n3537), .Y(n1898) );
  OAI21X1 U619 ( .A(n5771), .B(n5828), .C(n3614), .Y(n1899) );
  OAI21X1 U621 ( .A(n5772), .B(n5828), .C(n3075), .Y(n1900) );
  OAI21X1 U623 ( .A(n5748), .B(n5828), .C(n3459), .Y(n1901) );
  OAI21X1 U625 ( .A(n5747), .B(n5828), .C(n167), .Y(n1902) );
  OAI21X1 U628 ( .A(n5746), .B(n5827), .C(n3775), .Y(n1903) );
  OAI21X1 U630 ( .A(n5745), .B(n5826), .C(n3693), .Y(n1904) );
  OAI21X1 U632 ( .A(n5744), .B(n5827), .C(n3939), .Y(n1905) );
  OAI21X1 U634 ( .A(n5743), .B(n5827), .C(n3857), .Y(n1906) );
  OAI21X1 U636 ( .A(n5742), .B(n5827), .C(n4121), .Y(n1907) );
  OAI21X1 U638 ( .A(n5741), .B(n5826), .C(n4032), .Y(n1908) );
  OAI21X1 U640 ( .A(n5740), .B(n5826), .C(n4301), .Y(n1909) );
  OAI21X1 U642 ( .A(n5739), .B(n5826), .C(n4210), .Y(n1910) );
  OAI21X1 U644 ( .A(n5738), .B(n5827), .C(n3774), .Y(n1911) );
  OAI21X1 U646 ( .A(n5737), .B(n5826), .C(n3151), .Y(n1912) );
  OAI21X1 U648 ( .A(n5736), .B(n5826), .C(n3074), .Y(n1913) );
  OAI21X1 U650 ( .A(n5735), .B(n5827), .C(n3304), .Y(n1914) );
  OAI21X1 U652 ( .A(n5734), .B(n5826), .C(n3228), .Y(n1915) );
  OAI21X1 U654 ( .A(n5733), .B(n5826), .C(n3692), .Y(n1916) );
  OAI21X1 U656 ( .A(n5732), .B(n5827), .C(n3938), .Y(n1917) );
  OAI21X1 U658 ( .A(n5731), .B(n5826), .C(n3856), .Y(n1918) );
  OAI21X1 U660 ( .A(n5749), .B(n5827), .C(n3150), .Y(n1919) );
  OAI21X1 U662 ( .A(n5750), .B(n5826), .C(n4120), .Y(n1920) );
  OAI21X1 U664 ( .A(n5751), .B(n5827), .C(n4031), .Y(n1921) );
  OAI21X1 U666 ( .A(n5752), .B(n5826), .C(n4300), .Y(n1922) );
  OAI21X1 U668 ( .A(n5753), .B(n5827), .C(n4209), .Y(n1923) );
  OAI21X1 U670 ( .A(n5754), .B(n5826), .C(n3773), .Y(n1924) );
  OAI21X1 U672 ( .A(n5755), .B(n5826), .C(n3073), .Y(n1925) );
  OAI21X1 U674 ( .A(n5756), .B(n5827), .C(n3303), .Y(n1926) );
  OAI21X1 U676 ( .A(n5757), .B(n5827), .C(n3227), .Y(n1927) );
  OAI21X1 U678 ( .A(n5758), .B(n5827), .C(n3691), .Y(n1928) );
  OAI21X1 U680 ( .A(n5759), .B(n5827), .C(n3937), .Y(n1929) );
  OAI21X1 U682 ( .A(n5760), .B(n5826), .C(n4030), .Y(n1930) );
  OAI21X1 U684 ( .A(n5761), .B(n5826), .C(n4299), .Y(n1931) );
  OAI21X1 U686 ( .A(n5762), .B(n5827), .C(n4208), .Y(n1932) );
  OAI21X1 U688 ( .A(n5763), .B(n5827), .C(n3226), .Y(n1933) );
  OAI21X1 U690 ( .A(n5764), .B(n5826), .C(n3458), .Y(n1934) );
  OAI21X1 U692 ( .A(n5765), .B(n5826), .C(n3380), .Y(n1935) );
  OAI21X1 U694 ( .A(n5766), .B(n5826), .C(n3613), .Y(n1936) );
  OAI21X1 U696 ( .A(n5767), .B(n5827), .C(n3536), .Y(n1937) );
  OAI21X1 U698 ( .A(n5768), .B(n5826), .C(n166), .Y(n1938) );
  OAI21X1 U700 ( .A(n5769), .B(n5827), .C(n3072), .Y(n1939) );
  OAI21X1 U702 ( .A(n5770), .B(n5826), .C(n3457), .Y(n1940) );
  OAI21X1 U704 ( .A(n5771), .B(n5826), .C(n3379), .Y(n1941) );
  OAI21X1 U706 ( .A(n5772), .B(n5826), .C(n3302), .Y(n1942) );
  OAI21X1 U708 ( .A(n5748), .B(n5826), .C(n3535), .Y(n1943) );
  OAI21X1 U710 ( .A(n5747), .B(n5826), .C(n165), .Y(n1944) );
  OAI21X1 U713 ( .A(n5746), .B(n5825), .C(n3690), .Y(n1945) );
  OAI21X1 U715 ( .A(n5745), .B(n5824), .C(n3772), .Y(n1946) );
  OAI21X1 U717 ( .A(n5744), .B(n5825), .C(n3855), .Y(n1947) );
  OAI21X1 U719 ( .A(n5743), .B(n5825), .C(n3936), .Y(n1948) );
  OAI21X1 U721 ( .A(n5742), .B(n5825), .C(n4029), .Y(n1949) );
  OAI21X1 U723 ( .A(n5741), .B(n5824), .C(n4119), .Y(n1950) );
  OAI21X1 U725 ( .A(n5740), .B(n5824), .C(n4207), .Y(n1951) );
  OAI21X1 U727 ( .A(n5739), .B(n5824), .C(n4298), .Y(n1952) );
  OAI21X1 U729 ( .A(n5738), .B(n5825), .C(n3689), .Y(n1953) );
  OAI21X1 U731 ( .A(n5737), .B(n5824), .C(n3071), .Y(n1954) );
  OAI21X1 U733 ( .A(n5736), .B(n5824), .C(n3149), .Y(n1955) );
  OAI21X1 U735 ( .A(n5735), .B(n5825), .C(n3225), .Y(n1956) );
  OAI21X1 U737 ( .A(n5734), .B(n5824), .C(n3301), .Y(n1957) );
  OAI21X1 U739 ( .A(n5733), .B(n5824), .C(n3771), .Y(n1958) );
  OAI21X1 U741 ( .A(n5732), .B(n5825), .C(n3854), .Y(n1959) );
  OAI21X1 U743 ( .A(n5731), .B(n5824), .C(n3935), .Y(n1960) );
  OAI21X1 U745 ( .A(n5749), .B(n5825), .C(n3070), .Y(n1961) );
  OAI21X1 U747 ( .A(n5750), .B(n5824), .C(n4028), .Y(n1962) );
  OAI21X1 U749 ( .A(n5751), .B(n5825), .C(n4118), .Y(n1963) );
  OAI21X1 U751 ( .A(n5752), .B(n5824), .C(n4206), .Y(n1964) );
  OAI21X1 U753 ( .A(n5753), .B(n5825), .C(n4297), .Y(n1965) );
  OAI21X1 U755 ( .A(n5754), .B(n5824), .C(n3688), .Y(n1966) );
  OAI21X1 U757 ( .A(n5755), .B(n5824), .C(n3148), .Y(n1967) );
  OAI21X1 U759 ( .A(n5756), .B(n5825), .C(n3224), .Y(n1968) );
  OAI21X1 U761 ( .A(n5757), .B(n5825), .C(n3300), .Y(n1969) );
  OAI21X1 U763 ( .A(n5758), .B(n5825), .C(n3770), .Y(n1970) );
  OAI21X1 U765 ( .A(n5759), .B(n5825), .C(n3853), .Y(n1971) );
  OAI21X1 U767 ( .A(n5760), .B(n5824), .C(n4117), .Y(n1972) );
  OAI21X1 U769 ( .A(n5761), .B(n5824), .C(n4205), .Y(n1973) );
  OAI21X1 U771 ( .A(n5762), .B(n5825), .C(n4296), .Y(n1974) );
  OAI21X1 U773 ( .A(n5763), .B(n5825), .C(n3299), .Y(n1975) );
  OAI21X1 U775 ( .A(n5764), .B(n5824), .C(n3378), .Y(n1976) );
  OAI21X1 U777 ( .A(n5765), .B(n5824), .C(n3456), .Y(n1977) );
  OAI21X1 U779 ( .A(n5766), .B(n5824), .C(n3534), .Y(n1978) );
  OAI21X1 U781 ( .A(n5767), .B(n5825), .C(n3612), .Y(n1979) );
  OAI21X1 U783 ( .A(n5768), .B(n5824), .C(n164), .Y(n1980) );
  OAI21X1 U785 ( .A(n5769), .B(n5825), .C(n3147), .Y(n1981) );
  OAI21X1 U787 ( .A(n5770), .B(n5824), .C(n3377), .Y(n1982) );
  OAI21X1 U789 ( .A(n5771), .B(n5824), .C(n3455), .Y(n1983) );
  OAI21X1 U791 ( .A(n5772), .B(n5824), .C(n3223), .Y(n1984) );
  OAI21X1 U793 ( .A(n5748), .B(n5824), .C(n3611), .Y(n1985) );
  OAI21X1 U795 ( .A(n5747), .B(n5824), .C(n163), .Y(n1986) );
  NOR3X1 U798 ( .A(wr_ptr[3]), .B(wr_ptr[4]), .C(n1568), .Y(n222) );
  OAI21X1 U799 ( .A(n5746), .B(n5823), .C(n3610), .Y(n1987) );
  OAI21X1 U801 ( .A(n5745), .B(n5822), .C(n3533), .Y(n1988) );
  OAI21X1 U803 ( .A(n5744), .B(n5823), .C(n3454), .Y(n1989) );
  OAI21X1 U805 ( .A(n5743), .B(n5823), .C(n3376), .Y(n1990) );
  OAI21X1 U807 ( .A(n5742), .B(n5823), .C(n3298), .Y(n1991) );
  OAI21X1 U809 ( .A(n5741), .B(n5822), .C(n3222), .Y(n1992) );
  OAI21X1 U811 ( .A(n5740), .B(n5822), .C(n3146), .Y(n1993) );
  OAI21X1 U813 ( .A(n5739), .B(n5822), .C(n3069), .Y(n1994) );
  OAI21X1 U815 ( .A(n5738), .B(n5823), .C(n3609), .Y(n1995) );
  OAI21X1 U817 ( .A(n5737), .B(n5822), .C(n4295), .Y(n1996) );
  OAI21X1 U819 ( .A(n5736), .B(n5822), .C(n4204), .Y(n1997) );
  OAI21X1 U821 ( .A(n5735), .B(n5823), .C(n4116), .Y(n1998) );
  OAI21X1 U823 ( .A(n5734), .B(n5822), .C(n4027), .Y(n1999) );
  OAI21X1 U825 ( .A(n5733), .B(n5822), .C(n3532), .Y(n2000) );
  OAI21X1 U827 ( .A(n5732), .B(n5823), .C(n3453), .Y(n2001) );
  OAI21X1 U829 ( .A(n5731), .B(n5822), .C(n3375), .Y(n2002) );
  OAI21X1 U831 ( .A(n5749), .B(n5823), .C(n4294), .Y(n2003) );
  OAI21X1 U833 ( .A(n5750), .B(n5822), .C(n3297), .Y(n2004) );
  OAI21X1 U835 ( .A(n5751), .B(n5823), .C(n3221), .Y(n2005) );
  OAI21X1 U837 ( .A(n5752), .B(n5822), .C(n3145), .Y(n2006) );
  OAI21X1 U839 ( .A(n5753), .B(n5823), .C(n3068), .Y(n2007) );
  OAI21X1 U841 ( .A(n5754), .B(n5822), .C(n3608), .Y(n2008) );
  OAI21X1 U843 ( .A(n5755), .B(n5822), .C(n4203), .Y(n2009) );
  OAI21X1 U845 ( .A(n5756), .B(n5823), .C(n4115), .Y(n2010) );
  OAI21X1 U847 ( .A(n5757), .B(n5823), .C(n4026), .Y(n2011) );
  OAI21X1 U849 ( .A(n5758), .B(n5823), .C(n3531), .Y(n2012) );
  OAI21X1 U851 ( .A(n5759), .B(n5823), .C(n3452), .Y(n2013) );
  OAI21X1 U853 ( .A(n5760), .B(n5822), .C(n3220), .Y(n2014) );
  OAI21X1 U855 ( .A(n5761), .B(n5822), .C(n3144), .Y(n2015) );
  OAI21X1 U857 ( .A(n5762), .B(n5823), .C(n3067), .Y(n2016) );
  OAI21X1 U859 ( .A(n5763), .B(n5823), .C(n4025), .Y(n2017) );
  OAI21X1 U861 ( .A(n5764), .B(n5822), .C(n3934), .Y(n2018) );
  OAI21X1 U863 ( .A(n5765), .B(n5822), .C(n3852), .Y(n2019) );
  OAI21X1 U865 ( .A(n5766), .B(n5822), .C(n3769), .Y(n2020) );
  OAI21X1 U867 ( .A(n5767), .B(n5823), .C(n3687), .Y(n2021) );
  OAI21X1 U869 ( .A(n5768), .B(n5822), .C(n162), .Y(n2022) );
  OAI21X1 U871 ( .A(n5769), .B(n5823), .C(n4202), .Y(n2023) );
  OAI21X1 U873 ( .A(n5770), .B(n5822), .C(n3933), .Y(n2024) );
  OAI21X1 U875 ( .A(n5771), .B(n5822), .C(n3851), .Y(n2025) );
  OAI21X1 U877 ( .A(n5772), .B(n5822), .C(n4114), .Y(n2026) );
  OAI21X1 U879 ( .A(n5748), .B(n5822), .C(n3686), .Y(n2027) );
  OAI21X1 U881 ( .A(n5747), .B(n5822), .C(n161), .Y(n2028) );
  OAI21X1 U884 ( .A(n5746), .B(n5821), .C(n3530), .Y(n2029) );
  OAI21X1 U886 ( .A(n5745), .B(n5820), .C(n3607), .Y(n2030) );
  OAI21X1 U888 ( .A(n5744), .B(n5821), .C(n3374), .Y(n2031) );
  OAI21X1 U890 ( .A(n5743), .B(n5821), .C(n3451), .Y(n2032) );
  OAI21X1 U892 ( .A(n5742), .B(n5821), .C(n3219), .Y(n2033) );
  OAI21X1 U894 ( .A(n5741), .B(n5820), .C(n3296), .Y(n2034) );
  OAI21X1 U896 ( .A(n5740), .B(n5820), .C(n3066), .Y(n2035) );
  OAI21X1 U898 ( .A(n5739), .B(n5820), .C(n3143), .Y(n2036) );
  OAI21X1 U900 ( .A(n5738), .B(n5821), .C(n3529), .Y(n2037) );
  OAI21X1 U902 ( .A(n5737), .B(n5820), .C(n4201), .Y(n2038) );
  OAI21X1 U904 ( .A(n5736), .B(n5820), .C(n4293), .Y(n2039) );
  OAI21X1 U906 ( .A(n5735), .B(n5821), .C(n4024), .Y(n2040) );
  OAI21X1 U908 ( .A(n5734), .B(n5820), .C(n4113), .Y(n2041) );
  OAI21X1 U910 ( .A(n5733), .B(n5820), .C(n3606), .Y(n2042) );
  OAI21X1 U912 ( .A(n5732), .B(n5821), .C(n3373), .Y(n2043) );
  OAI21X1 U914 ( .A(n5731), .B(n5820), .C(n3450), .Y(n2044) );
  OAI21X1 U916 ( .A(n5749), .B(n5821), .C(n4200), .Y(n2045) );
  OAI21X1 U918 ( .A(n5750), .B(n5820), .C(n3218), .Y(n2046) );
  OAI21X1 U920 ( .A(n5751), .B(n5821), .C(n3295), .Y(n2047) );
  OAI21X1 U922 ( .A(n5752), .B(n5820), .C(n3065), .Y(n2048) );
  OAI21X1 U924 ( .A(n5753), .B(n5821), .C(n3142), .Y(n2049) );
  OAI21X1 U926 ( .A(n5754), .B(n5820), .C(n3528), .Y(n2050) );
  OAI21X1 U928 ( .A(n5755), .B(n5820), .C(n4292), .Y(n2051) );
  OAI21X1 U930 ( .A(n5756), .B(n5821), .C(n4023), .Y(n2052) );
  OAI21X1 U932 ( .A(n5757), .B(n5821), .C(n4112), .Y(n2053) );
  OAI21X1 U934 ( .A(n5758), .B(n5821), .C(n3605), .Y(n2054) );
  OAI21X1 U936 ( .A(n5759), .B(n5821), .C(n3372), .Y(n2055) );
  OAI21X1 U938 ( .A(n5760), .B(n5820), .C(n3294), .Y(n2056) );
  OAI21X1 U940 ( .A(n5761), .B(n5820), .C(n3064), .Y(n2057) );
  OAI21X1 U942 ( .A(n5762), .B(n5821), .C(n3141), .Y(n2058) );
  OAI21X1 U944 ( .A(n5763), .B(n5821), .C(n4111), .Y(n2059) );
  OAI21X1 U946 ( .A(n5764), .B(n5820), .C(n3850), .Y(n2060) );
  OAI21X1 U948 ( .A(n5765), .B(n5820), .C(n3932), .Y(n2061) );
  OAI21X1 U950 ( .A(n5766), .B(n5820), .C(n3685), .Y(n2062) );
  OAI21X1 U952 ( .A(n5767), .B(n5821), .C(n3768), .Y(n2063) );
  OAI21X1 U954 ( .A(n5768), .B(n5820), .C(n160), .Y(n2064) );
  OAI21X1 U956 ( .A(n5769), .B(n5821), .C(n4291), .Y(n2065) );
  OAI21X1 U958 ( .A(n5770), .B(n5820), .C(n3849), .Y(n2066) );
  OAI21X1 U960 ( .A(n5771), .B(n5820), .C(n3931), .Y(n2067) );
  OAI21X1 U962 ( .A(n5772), .B(n5820), .C(n4022), .Y(n2068) );
  OAI21X1 U964 ( .A(n5748), .B(n5820), .C(n3767), .Y(n2069) );
  OAI21X1 U966 ( .A(n5747), .B(n5820), .C(n159), .Y(n2070) );
  OAI21X1 U969 ( .A(n5746), .B(n5819), .C(n3449), .Y(n2071) );
  OAI21X1 U971 ( .A(n5745), .B(n5818), .C(n3371), .Y(n2072) );
  OAI21X1 U973 ( .A(n5744), .B(n5819), .C(n3604), .Y(n2073) );
  OAI21X1 U975 ( .A(n5743), .B(n5819), .C(n3527), .Y(n2074) );
  OAI21X1 U977 ( .A(n5742), .B(n5819), .C(n3140), .Y(n2075) );
  OAI21X1 U979 ( .A(n5741), .B(n5818), .C(n3063), .Y(n2076) );
  OAI21X1 U981 ( .A(n5740), .B(n5818), .C(n3293), .Y(n2077) );
  OAI21X1 U983 ( .A(n5739), .B(n5818), .C(n3217), .Y(n2078) );
  OAI21X1 U985 ( .A(n5738), .B(n5819), .C(n3448), .Y(n2079) );
  OAI21X1 U987 ( .A(n5737), .B(n5818), .C(n4110), .Y(n2080) );
  OAI21X1 U989 ( .A(n5736), .B(n5818), .C(n4021), .Y(n2081) );
  OAI21X1 U991 ( .A(n5735), .B(n5819), .C(n4290), .Y(n2082) );
  OAI21X1 U993 ( .A(n5734), .B(n5818), .C(n4199), .Y(n2083) );
  OAI21X1 U995 ( .A(n5733), .B(n5818), .C(n3370), .Y(n2084) );
  OAI21X1 U997 ( .A(n5732), .B(n5819), .C(n3603), .Y(n2085) );
  OAI21X1 U999 ( .A(n5731), .B(n5818), .C(n3526), .Y(n2086) );
  OAI21X1 U1001 ( .A(n5749), .B(n5819), .C(n4109), .Y(n2087) );
  OAI21X1 U1003 ( .A(n5750), .B(n5818), .C(n3139), .Y(n2088) );
  OAI21X1 U1005 ( .A(n5751), .B(n5819), .C(n3062), .Y(n2089) );
  OAI21X1 U1007 ( .A(n5752), .B(n5818), .C(n3292), .Y(n2090) );
  OAI21X1 U1009 ( .A(n5753), .B(n5819), .C(n3216), .Y(n2091) );
  OAI21X1 U1011 ( .A(n5754), .B(n5818), .C(n3447), .Y(n2092) );
  OAI21X1 U1013 ( .A(n5755), .B(n5818), .C(n4020), .Y(n2093) );
  OAI21X1 U1015 ( .A(n5756), .B(n5819), .C(n4289), .Y(n2094) );
  OAI21X1 U1017 ( .A(n5757), .B(n5819), .C(n4198), .Y(n2095) );
  OAI21X1 U1019 ( .A(n5758), .B(n5819), .C(n3369), .Y(n2096) );
  OAI21X1 U1021 ( .A(n5759), .B(n5819), .C(n3602), .Y(n2097) );
  OAI21X1 U1023 ( .A(n5760), .B(n5818), .C(n3061), .Y(n2098) );
  OAI21X1 U1025 ( .A(n5761), .B(n5818), .C(n3291), .Y(n2099) );
  OAI21X1 U1027 ( .A(n5762), .B(n5819), .C(n3215), .Y(n2100) );
  OAI21X1 U1029 ( .A(n5763), .B(n5819), .C(n4197), .Y(n2101) );
  OAI21X1 U1031 ( .A(n5764), .B(n5818), .C(n3766), .Y(n2102) );
  OAI21X1 U1033 ( .A(n5765), .B(n5818), .C(n3684), .Y(n2103) );
  OAI21X1 U1035 ( .A(n5766), .B(n5818), .C(n3930), .Y(n2104) );
  OAI21X1 U1037 ( .A(n5767), .B(n5819), .C(n3848), .Y(n2105) );
  OAI21X1 U1039 ( .A(n5768), .B(n5818), .C(n158), .Y(n2106) );
  OAI21X1 U1041 ( .A(n5769), .B(n5819), .C(n4019), .Y(n2107) );
  OAI21X1 U1043 ( .A(n5770), .B(n5818), .C(n3765), .Y(n2108) );
  OAI21X1 U1045 ( .A(n5771), .B(n5818), .C(n3683), .Y(n2109) );
  OAI21X1 U1047 ( .A(n5772), .B(n5818), .C(n4288), .Y(n2110) );
  OAI21X1 U1049 ( .A(n5748), .B(n5818), .C(n3847), .Y(n2111) );
  OAI21X1 U1051 ( .A(n5747), .B(n5818), .C(n157), .Y(n2112) );
  OAI21X1 U1054 ( .A(n5746), .B(n5817), .C(n3368), .Y(n2113) );
  OAI21X1 U1056 ( .A(n5745), .B(n5816), .C(n3446), .Y(n2114) );
  OAI21X1 U1058 ( .A(n5744), .B(n5817), .C(n3525), .Y(n2115) );
  OAI21X1 U1060 ( .A(n5743), .B(n5817), .C(n3601), .Y(n2116) );
  OAI21X1 U1062 ( .A(n5742), .B(n5817), .C(n3060), .Y(n2117) );
  OAI21X1 U1064 ( .A(n5741), .B(n5816), .C(n3138), .Y(n2118) );
  OAI21X1 U1066 ( .A(n5740), .B(n5816), .C(n3214), .Y(n2119) );
  OAI21X1 U1068 ( .A(n5739), .B(n5816), .C(n3290), .Y(n2120) );
  OAI21X1 U1070 ( .A(n5738), .B(n5817), .C(n3367), .Y(n2121) );
  OAI21X1 U1072 ( .A(n5737), .B(n5816), .C(n4018), .Y(n2122) );
  OAI21X1 U1074 ( .A(n5736), .B(n5816), .C(n4108), .Y(n2123) );
  OAI21X1 U1076 ( .A(n5735), .B(n5817), .C(n4196), .Y(n2124) );
  OAI21X1 U1078 ( .A(n5734), .B(n5816), .C(n4287), .Y(n2125) );
  OAI21X1 U1080 ( .A(n5733), .B(n5816), .C(n3445), .Y(n2126) );
  OAI21X1 U1082 ( .A(n5732), .B(n5817), .C(n3524), .Y(n2127) );
  OAI21X1 U1084 ( .A(n5731), .B(n5816), .C(n3600), .Y(n2128) );
  OAI21X1 U1086 ( .A(n5749), .B(n5817), .C(n4017), .Y(n2129) );
  OAI21X1 U1088 ( .A(n5750), .B(n5816), .C(n3059), .Y(n2130) );
  OAI21X1 U1090 ( .A(n5751), .B(n5817), .C(n3137), .Y(n2131) );
  OAI21X1 U1092 ( .A(n5752), .B(n5816), .C(n3213), .Y(n2132) );
  OAI21X1 U1094 ( .A(n5753), .B(n5817), .C(n3289), .Y(n2133) );
  OAI21X1 U1096 ( .A(n5754), .B(n5816), .C(n3366), .Y(n2134) );
  OAI21X1 U1098 ( .A(n5755), .B(n5816), .C(n4107), .Y(n2135) );
  OAI21X1 U1100 ( .A(n5756), .B(n5817), .C(n4195), .Y(n2136) );
  OAI21X1 U1102 ( .A(n5757), .B(n5817), .C(n4286), .Y(n2137) );
  OAI21X1 U1104 ( .A(n5758), .B(n5817), .C(n3444), .Y(n2138) );
  OAI21X1 U1106 ( .A(n5759), .B(n5817), .C(n3523), .Y(n2139) );
  OAI21X1 U1108 ( .A(n5760), .B(n5816), .C(n3136), .Y(n2140) );
  OAI21X1 U1110 ( .A(n5761), .B(n5816), .C(n3212), .Y(n2141) );
  OAI21X1 U1112 ( .A(n5762), .B(n5817), .C(n3288), .Y(n2142) );
  OAI21X1 U1114 ( .A(n5763), .B(n5817), .C(n4285), .Y(n2143) );
  OAI21X1 U1116 ( .A(n5764), .B(n5816), .C(n3682), .Y(n2144) );
  OAI21X1 U1118 ( .A(n5765), .B(n5816), .C(n3764), .Y(n2145) );
  OAI21X1 U1120 ( .A(n5766), .B(n5816), .C(n3846), .Y(n2146) );
  OAI21X1 U1122 ( .A(n5767), .B(n5817), .C(n3929), .Y(n2147) );
  OAI21X1 U1124 ( .A(n5768), .B(n5816), .C(n156), .Y(n2148) );
  OAI21X1 U1126 ( .A(n5769), .B(n5817), .C(n4106), .Y(n2149) );
  OAI21X1 U1128 ( .A(n5770), .B(n5816), .C(n3681), .Y(n2150) );
  OAI21X1 U1130 ( .A(n5771), .B(n5816), .C(n3763), .Y(n2151) );
  OAI21X1 U1132 ( .A(n5772), .B(n5816), .C(n4194), .Y(n2152) );
  OAI21X1 U1134 ( .A(n5748), .B(n5816), .C(n3928), .Y(n2153) );
  OAI21X1 U1136 ( .A(n5747), .B(n5816), .C(n155), .Y(n2154) );
  OAI21X1 U1139 ( .A(n5746), .B(n5815), .C(n3287), .Y(n2155) );
  OAI21X1 U1141 ( .A(n5745), .B(n5814), .C(n3211), .Y(n2156) );
  OAI21X1 U1143 ( .A(n5744), .B(n5815), .C(n3135), .Y(n2157) );
  OAI21X1 U1145 ( .A(n5743), .B(n5815), .C(n3058), .Y(n2158) );
  OAI21X1 U1147 ( .A(n5742), .B(n5815), .C(n3599), .Y(n2159) );
  OAI21X1 U1149 ( .A(n5741), .B(n5814), .C(n3522), .Y(n2160) );
  OAI21X1 U1151 ( .A(n5740), .B(n5814), .C(n3443), .Y(n2161) );
  OAI21X1 U1153 ( .A(n5739), .B(n5814), .C(n3365), .Y(n2162) );
  OAI21X1 U1155 ( .A(n5738), .B(n5815), .C(n3286), .Y(n2163) );
  OAI21X1 U1157 ( .A(n5737), .B(n5814), .C(n3927), .Y(n2164) );
  OAI21X1 U1159 ( .A(n5736), .B(n5814), .C(n3845), .Y(n2165) );
  OAI21X1 U1161 ( .A(n5735), .B(n5815), .C(n3762), .Y(n2166) );
  OAI21X1 U1163 ( .A(n5734), .B(n5814), .C(n3680), .Y(n2167) );
  OAI21X1 U1165 ( .A(n5733), .B(n5814), .C(n3210), .Y(n2168) );
  OAI21X1 U1167 ( .A(n5732), .B(n5815), .C(n3134), .Y(n2169) );
  OAI21X1 U1169 ( .A(n5731), .B(n5814), .C(n3057), .Y(n2170) );
  OAI21X1 U1171 ( .A(n5749), .B(n5815), .C(n3926), .Y(n2171) );
  OAI21X1 U1173 ( .A(n5750), .B(n5814), .C(n3598), .Y(n2172) );
  OAI21X1 U1175 ( .A(n5751), .B(n5815), .C(n3521), .Y(n2173) );
  OAI21X1 U1177 ( .A(n5752), .B(n5814), .C(n3442), .Y(n2174) );
  OAI21X1 U1179 ( .A(n5753), .B(n5815), .C(n3364), .Y(n2175) );
  OAI21X1 U1181 ( .A(n5754), .B(n5814), .C(n3285), .Y(n2176) );
  OAI21X1 U1183 ( .A(n5755), .B(n5814), .C(n3844), .Y(n2177) );
  OAI21X1 U1185 ( .A(n5756), .B(n5815), .C(n3761), .Y(n2178) );
  OAI21X1 U1187 ( .A(n5757), .B(n5815), .C(n3679), .Y(n2179) );
  OAI21X1 U1189 ( .A(n5758), .B(n5815), .C(n3209), .Y(n2180) );
  OAI21X1 U1191 ( .A(n5759), .B(n5815), .C(n3133), .Y(n2181) );
  OAI21X1 U1193 ( .A(n5760), .B(n5814), .C(n3520), .Y(n2182) );
  OAI21X1 U1195 ( .A(n5761), .B(n5814), .C(n3441), .Y(n2183) );
  OAI21X1 U1197 ( .A(n5762), .B(n5815), .C(n3363), .Y(n2184) );
  OAI21X1 U1199 ( .A(n5763), .B(n5815), .C(n3678), .Y(n2185) );
  OAI21X1 U1201 ( .A(n5764), .B(n5814), .C(n4284), .Y(n2186) );
  OAI21X1 U1203 ( .A(n5765), .B(n5814), .C(n4193), .Y(n2187) );
  OAI21X1 U1205 ( .A(n5766), .B(n5814), .C(n4105), .Y(n2188) );
  OAI21X1 U1207 ( .A(n5767), .B(n5815), .C(n4016), .Y(n2189) );
  OAI21X1 U1209 ( .A(n5768), .B(n5814), .C(n154), .Y(n2190) );
  OAI21X1 U1211 ( .A(n5769), .B(n5815), .C(n3843), .Y(n2191) );
  OAI21X1 U1213 ( .A(n5770), .B(n5814), .C(n4283), .Y(n2192) );
  OAI21X1 U1215 ( .A(n5771), .B(n5814), .C(n4192), .Y(n2193) );
  OAI21X1 U1217 ( .A(n5772), .B(n5814), .C(n3760), .Y(n2194) );
  OAI21X1 U1219 ( .A(n5748), .B(n5814), .C(n4015), .Y(n2195) );
  OAI21X1 U1221 ( .A(n5747), .B(n5814), .C(n153), .Y(n2196) );
  OAI21X1 U1224 ( .A(n5746), .B(n5812), .C(n4282), .Y(n2197) );
  OAI21X1 U1226 ( .A(n5745), .B(n5812), .C(n4191), .Y(n2198) );
  OAI21X1 U1228 ( .A(n5744), .B(n5812), .C(n4104), .Y(n2199) );
  OAI21X1 U1230 ( .A(n5743), .B(n5812), .C(n4014), .Y(n2200) );
  OAI21X1 U1232 ( .A(n5742), .B(n5813), .C(n3925), .Y(n2201) );
  OAI21X1 U1234 ( .A(n5741), .B(n5812), .C(n3842), .Y(n2202) );
  OAI21X1 U1236 ( .A(n5740), .B(n5813), .C(n3759), .Y(n2203) );
  OAI21X1 U1238 ( .A(n5739), .B(n5812), .C(n3677), .Y(n2204) );
  OAI21X1 U1240 ( .A(n5738), .B(n5813), .C(n4281), .Y(n2205) );
  OAI21X1 U1242 ( .A(n5737), .B(n5813), .C(n3597), .Y(n2206) );
  OAI21X1 U1244 ( .A(n5736), .B(n5813), .C(n3519), .Y(n2207) );
  OAI21X1 U1246 ( .A(n5735), .B(n5813), .C(n3440), .Y(n2208) );
  OAI21X1 U1248 ( .A(n5734), .B(n5812), .C(n3362), .Y(n2209) );
  OAI21X1 U1250 ( .A(n5733), .B(n5812), .C(n4190), .Y(n2210) );
  OAI21X1 U1252 ( .A(n5732), .B(n5812), .C(n4103), .Y(n2211) );
  OAI21X1 U1254 ( .A(n5731), .B(n5813), .C(n4013), .Y(n2212) );
  OAI21X1 U1256 ( .A(n5749), .B(n5813), .C(n3596), .Y(n2213) );
  OAI21X1 U1258 ( .A(n5750), .B(n5812), .C(n3924), .Y(n2214) );
  OAI21X1 U1260 ( .A(n5751), .B(n5813), .C(n3841), .Y(n2215) );
  OAI21X1 U1262 ( .A(n5752), .B(n5813), .C(n3758), .Y(n2216) );
  OAI21X1 U1264 ( .A(n5753), .B(n5813), .C(n3676), .Y(n2217) );
  OAI21X1 U1266 ( .A(n5754), .B(n5813), .C(n4280), .Y(n2218) );
  OAI21X1 U1268 ( .A(n5755), .B(n5812), .C(n3518), .Y(n2219) );
  OAI21X1 U1270 ( .A(n5756), .B(n5812), .C(n3439), .Y(n2220) );
  OAI21X1 U1272 ( .A(n5757), .B(n5813), .C(n3361), .Y(n2221) );
  OAI21X1 U1274 ( .A(n5758), .B(n5813), .C(n4189), .Y(n2222) );
  OAI21X1 U1276 ( .A(n5759), .B(n5812), .C(n4102), .Y(n2223) );
  OAI21X1 U1278 ( .A(n5760), .B(n5813), .C(n3840), .Y(n2224) );
  OAI21X1 U1280 ( .A(n5761), .B(n5812), .C(n3757), .Y(n2225) );
  OAI21X1 U1282 ( .A(n5762), .B(n5813), .C(n3675), .Y(n2226) );
  OAI21X1 U1284 ( .A(n5763), .B(n5812), .C(n3360), .Y(n2227) );
  OAI21X1 U1286 ( .A(n5764), .B(n5813), .C(n3284), .Y(n2228) );
  OAI21X1 U1288 ( .A(n5765), .B(n5812), .C(n3208), .Y(n2229) );
  OAI21X1 U1290 ( .A(n5766), .B(n5812), .C(n3132), .Y(n2230) );
  OAI21X1 U1292 ( .A(n5767), .B(n5812), .C(n3056), .Y(n2231) );
  OAI21X1 U1294 ( .A(n5768), .B(n5812), .C(n152), .Y(n2232) );
  OAI21X1 U1296 ( .A(n5769), .B(n5812), .C(n3517), .Y(n2233) );
  OAI21X1 U1298 ( .A(n5770), .B(n5812), .C(n3283), .Y(n2234) );
  OAI21X1 U1300 ( .A(n5771), .B(n5812), .C(n3207), .Y(n2235) );
  OAI21X1 U1302 ( .A(n5772), .B(n5813), .C(n3438), .Y(n2236) );
  OAI21X1 U1304 ( .A(n5748), .B(n5812), .C(n3055), .Y(n2237) );
  OAI21X1 U1306 ( .A(n5747), .B(n5812), .C(n151), .Y(n2238) );
  OAI21X1 U1309 ( .A(n5746), .B(n5810), .C(n4188), .Y(n2239) );
  OAI21X1 U1311 ( .A(n5745), .B(n5810), .C(n4279), .Y(n2240) );
  OAI21X1 U1313 ( .A(n5744), .B(n5810), .C(n4012), .Y(n2241) );
  OAI21X1 U1315 ( .A(n5743), .B(n5810), .C(n4101), .Y(n2242) );
  OAI21X1 U1317 ( .A(n5742), .B(n5811), .C(n3839), .Y(n2243) );
  OAI21X1 U1319 ( .A(n5741), .B(n5810), .C(n3923), .Y(n2244) );
  OAI21X1 U1321 ( .A(n5740), .B(n5811), .C(n3674), .Y(n2245) );
  OAI21X1 U1323 ( .A(n5739), .B(n5810), .C(n3756), .Y(n2246) );
  OAI21X1 U1325 ( .A(n5738), .B(n5811), .C(n4187), .Y(n2247) );
  OAI21X1 U1327 ( .A(n5737), .B(n5811), .C(n3516), .Y(n2248) );
  OAI21X1 U1329 ( .A(n5736), .B(n5811), .C(n3595), .Y(n2249) );
  OAI21X1 U1331 ( .A(n5735), .B(n5811), .C(n3359), .Y(n2250) );
  OAI21X1 U1333 ( .A(n5734), .B(n5810), .C(n3437), .Y(n2251) );
  OAI21X1 U1335 ( .A(n5733), .B(n5810), .C(n4278), .Y(n2252) );
  OAI21X1 U1337 ( .A(n5732), .B(n5810), .C(n4011), .Y(n2253) );
  OAI21X1 U1339 ( .A(n5731), .B(n5811), .C(n4100), .Y(n2254) );
  OAI21X1 U1341 ( .A(n5749), .B(n5811), .C(n3515), .Y(n2255) );
  OAI21X1 U1343 ( .A(n5750), .B(n5810), .C(n3838), .Y(n2256) );
  OAI21X1 U1345 ( .A(n5751), .B(n5811), .C(n3922), .Y(n2257) );
  OAI21X1 U1347 ( .A(n5752), .B(n5811), .C(n3673), .Y(n2258) );
  OAI21X1 U1349 ( .A(n5753), .B(n5811), .C(n3755), .Y(n2259) );
  OAI21X1 U1351 ( .A(n5754), .B(n5811), .C(n4186), .Y(n2260) );
  OAI21X1 U1353 ( .A(n5755), .B(n5810), .C(n3594), .Y(n2261) );
  OAI21X1 U1355 ( .A(n5756), .B(n5810), .C(n3358), .Y(n2262) );
  OAI21X1 U1357 ( .A(n5757), .B(n5811), .C(n3436), .Y(n2263) );
  OAI21X1 U1359 ( .A(n5758), .B(n5811), .C(n4277), .Y(n2264) );
  OAI21X1 U1361 ( .A(n5759), .B(n5810), .C(n4010), .Y(n2265) );
  OAI21X1 U1363 ( .A(n5760), .B(n5811), .C(n3921), .Y(n2266) );
  OAI21X1 U1365 ( .A(n5761), .B(n5810), .C(n3672), .Y(n2267) );
  OAI21X1 U1367 ( .A(n5762), .B(n5811), .C(n3754), .Y(n2268) );
  OAI21X1 U1369 ( .A(n5763), .B(n5810), .C(n3435), .Y(n2269) );
  OAI21X1 U1371 ( .A(n5764), .B(n5811), .C(n3206), .Y(n2270) );
  OAI21X1 U1373 ( .A(n5765), .B(n5810), .C(n3282), .Y(n2271) );
  OAI21X1 U1375 ( .A(n5766), .B(n5810), .C(n3054), .Y(n2272) );
  OAI21X1 U1377 ( .A(n5767), .B(n5810), .C(n3131), .Y(n2273) );
  OAI21X1 U1379 ( .A(n5768), .B(n5810), .C(n150), .Y(n2274) );
  OAI21X1 U1381 ( .A(n5769), .B(n5810), .C(n3593), .Y(n2275) );
  OAI21X1 U1383 ( .A(n5770), .B(n5810), .C(n3205), .Y(n2276) );
  OAI21X1 U1385 ( .A(n5771), .B(n5810), .C(n3281), .Y(n2277) );
  OAI21X1 U1387 ( .A(n5772), .B(n5811), .C(n3357), .Y(n2278) );
  OAI21X1 U1389 ( .A(n5748), .B(n5810), .C(n3130), .Y(n2279) );
  OAI21X1 U1391 ( .A(n5747), .B(n5810), .C(n149), .Y(n2280) );
  OAI21X1 U1394 ( .A(n5746), .B(n5808), .C(n4099), .Y(n2281) );
  OAI21X1 U1396 ( .A(n5745), .B(n5808), .C(n4009), .Y(n2282) );
  OAI21X1 U1398 ( .A(n5744), .B(n5808), .C(n4276), .Y(n2283) );
  OAI21X1 U1400 ( .A(n5743), .B(n5808), .C(n4185), .Y(n2284) );
  OAI21X1 U1402 ( .A(n5742), .B(n5809), .C(n3753), .Y(n2285) );
  OAI21X1 U1404 ( .A(n5741), .B(n5808), .C(n3671), .Y(n2286) );
  OAI21X1 U1406 ( .A(n5740), .B(n5809), .C(n3920), .Y(n2287) );
  OAI21X1 U1408 ( .A(n5739), .B(n5808), .C(n3837), .Y(n2288) );
  OAI21X1 U1410 ( .A(n5738), .B(n5809), .C(n4098), .Y(n2289) );
  OAI21X1 U1412 ( .A(n5737), .B(n5809), .C(n3434), .Y(n2290) );
  OAI21X1 U1414 ( .A(n5736), .B(n5809), .C(n3356), .Y(n2291) );
  OAI21X1 U1416 ( .A(n5735), .B(n5809), .C(n3592), .Y(n2292) );
  OAI21X1 U1418 ( .A(n5734), .B(n5808), .C(n3514), .Y(n2293) );
  OAI21X1 U1420 ( .A(n5733), .B(n5808), .C(n4008), .Y(n2294) );
  OAI21X1 U1422 ( .A(n5732), .B(n5808), .C(n4275), .Y(n2295) );
  OAI21X1 U1424 ( .A(n5731), .B(n5809), .C(n4184), .Y(n2296) );
  OAI21X1 U1426 ( .A(n5749), .B(n5809), .C(n3433), .Y(n2297) );
  OAI21X1 U1428 ( .A(n5750), .B(n5808), .C(n3752), .Y(n2298) );
  OAI21X1 U1430 ( .A(n5751), .B(n5809), .C(n3670), .Y(n2299) );
  OAI21X1 U1432 ( .A(n5752), .B(n5809), .C(n3919), .Y(n2300) );
  OAI21X1 U1434 ( .A(n5753), .B(n5809), .C(n3836), .Y(n2301) );
  OAI21X1 U1436 ( .A(n5754), .B(n5809), .C(n4097), .Y(n2302) );
  OAI21X1 U1438 ( .A(n5755), .B(n5808), .C(n3355), .Y(n2303) );
  OAI21X1 U1440 ( .A(n5756), .B(n5808), .C(n3591), .Y(n2304) );
  OAI21X1 U1442 ( .A(n5757), .B(n5809), .C(n3513), .Y(n2305) );
  OAI21X1 U1444 ( .A(n5758), .B(n5809), .C(n4007), .Y(n2306) );
  OAI21X1 U1446 ( .A(n5759), .B(n5808), .C(n4274), .Y(n2307) );
  OAI21X1 U1448 ( .A(n5760), .B(n5809), .C(n3669), .Y(n2308) );
  OAI21X1 U1450 ( .A(n5761), .B(n5808), .C(n3918), .Y(n2309) );
  OAI21X1 U1452 ( .A(n5762), .B(n5809), .C(n3835), .Y(n2310) );
  OAI21X1 U1454 ( .A(n5763), .B(n5808), .C(n3512), .Y(n2311) );
  OAI21X1 U1456 ( .A(n5764), .B(n5809), .C(n3129), .Y(n2312) );
  OAI21X1 U1458 ( .A(n5765), .B(n5808), .C(n3053), .Y(n2313) );
  OAI21X1 U1460 ( .A(n5766), .B(n5808), .C(n3280), .Y(n2314) );
  OAI21X1 U1462 ( .A(n5767), .B(n5808), .C(n3204), .Y(n2315) );
  OAI21X1 U1464 ( .A(n5768), .B(n5808), .C(n148), .Y(n2316) );
  OAI21X1 U1466 ( .A(n5769), .B(n5808), .C(n3354), .Y(n2317) );
  OAI21X1 U1468 ( .A(n5770), .B(n5808), .C(n3128), .Y(n2318) );
  OAI21X1 U1470 ( .A(n5771), .B(n5808), .C(n3052), .Y(n2319) );
  OAI21X1 U1472 ( .A(n5772), .B(n5809), .C(n3590), .Y(n2320) );
  OAI21X1 U1474 ( .A(n5748), .B(n5808), .C(n3203), .Y(n2321) );
  OAI21X1 U1476 ( .A(n5747), .B(n5808), .C(n147), .Y(n2322) );
  NOR3X1 U1479 ( .A(n1568), .B(wr_ptr[4]), .C(n5901), .Y(n574) );
  OAI21X1 U1480 ( .A(n5746), .B(n5806), .C(n4006), .Y(n2323) );
  OAI21X1 U1482 ( .A(n5745), .B(n5806), .C(n4096), .Y(n2324) );
  OAI21X1 U1484 ( .A(n5744), .B(n5806), .C(n4183), .Y(n2325) );
  OAI21X1 U1486 ( .A(n5743), .B(n5806), .C(n4273), .Y(n2326) );
  OAI21X1 U1488 ( .A(n5742), .B(n5807), .C(n3668), .Y(n2327) );
  OAI21X1 U1490 ( .A(n5741), .B(n5806), .C(n3751), .Y(n2328) );
  OAI21X1 U1492 ( .A(n5740), .B(n5807), .C(n3834), .Y(n2329) );
  OAI21X1 U1494 ( .A(n5739), .B(n5806), .C(n3917), .Y(n2330) );
  OAI21X1 U1496 ( .A(n5738), .B(n5807), .C(n4005), .Y(n2331) );
  OAI21X1 U1498 ( .A(n5737), .B(n5807), .C(n3353), .Y(n2332) );
  OAI21X1 U1500 ( .A(n5736), .B(n5807), .C(n3432), .Y(n2333) );
  OAI21X1 U1502 ( .A(n5735), .B(n5807), .C(n3511), .Y(n2334) );
  OAI21X1 U1504 ( .A(n5734), .B(n5806), .C(n3589), .Y(n2335) );
  OAI21X1 U1506 ( .A(n5733), .B(n5806), .C(n4095), .Y(n2336) );
  OAI21X1 U1508 ( .A(n5732), .B(n5806), .C(n4182), .Y(n2337) );
  OAI21X1 U1510 ( .A(n5731), .B(n5807), .C(n4272), .Y(n2338) );
  OAI21X1 U1512 ( .A(n5749), .B(n5807), .C(n3352), .Y(n2339) );
  OAI21X1 U1514 ( .A(n5750), .B(n5806), .C(n3667), .Y(n2340) );
  OAI21X1 U1516 ( .A(n5751), .B(n5807), .C(n3750), .Y(n2341) );
  OAI21X1 U1518 ( .A(n5752), .B(n5807), .C(n3833), .Y(n2342) );
  OAI21X1 U1520 ( .A(n5753), .B(n5807), .C(n3916), .Y(n2343) );
  OAI21X1 U1522 ( .A(n5754), .B(n5807), .C(n4004), .Y(n2344) );
  OAI21X1 U1524 ( .A(n5755), .B(n5806), .C(n3431), .Y(n2345) );
  OAI21X1 U1526 ( .A(n5756), .B(n5806), .C(n3510), .Y(n2346) );
  OAI21X1 U1528 ( .A(n5757), .B(n5807), .C(n3588), .Y(n2347) );
  OAI21X1 U1530 ( .A(n5758), .B(n5807), .C(n4094), .Y(n2348) );
  OAI21X1 U1532 ( .A(n5759), .B(n5806), .C(n4181), .Y(n2349) );
  OAI21X1 U1534 ( .A(n5760), .B(n5807), .C(n3749), .Y(n2350) );
  OAI21X1 U1536 ( .A(n5761), .B(n5806), .C(n3832), .Y(n2351) );
  OAI21X1 U1538 ( .A(n5762), .B(n5807), .C(n3915), .Y(n2352) );
  OAI21X1 U1540 ( .A(n5763), .B(n5806), .C(n3587), .Y(n2353) );
  OAI21X1 U1542 ( .A(n5764), .B(n5807), .C(n3051), .Y(n2354) );
  OAI21X1 U1544 ( .A(n5765), .B(n5806), .C(n3127), .Y(n2355) );
  OAI21X1 U1546 ( .A(n5766), .B(n5806), .C(n3202), .Y(n2356) );
  OAI21X1 U1548 ( .A(n5767), .B(n5806), .C(n3279), .Y(n2357) );
  OAI21X1 U1550 ( .A(n5768), .B(n5806), .C(n146), .Y(n2358) );
  OAI21X1 U1552 ( .A(n5769), .B(n5806), .C(n3430), .Y(n2359) );
  OAI21X1 U1554 ( .A(n5770), .B(n5806), .C(n3050), .Y(n2360) );
  OAI21X1 U1556 ( .A(n5771), .B(n5806), .C(n3126), .Y(n2361) );
  OAI21X1 U1558 ( .A(n5772), .B(n5807), .C(n3509), .Y(n2362) );
  OAI21X1 U1560 ( .A(n5748), .B(n5806), .C(n3278), .Y(n2363) );
  OAI21X1 U1562 ( .A(n5747), .B(n5806), .C(n145), .Y(n2364) );
  OAI21X1 U1565 ( .A(n5746), .B(n5804), .C(n3914), .Y(n2365) );
  OAI21X1 U1567 ( .A(n5745), .B(n5804), .C(n3831), .Y(n2366) );
  OAI21X1 U1569 ( .A(n5744), .B(n5804), .C(n3748), .Y(n2367) );
  OAI21X1 U1571 ( .A(n5743), .B(n5804), .C(n3666), .Y(n2368) );
  OAI21X1 U1573 ( .A(n5742), .B(n5805), .C(n4271), .Y(n2369) );
  OAI21X1 U1575 ( .A(n5741), .B(n5804), .C(n4180), .Y(n2370) );
  OAI21X1 U1577 ( .A(n5740), .B(n5805), .C(n4093), .Y(n2371) );
  OAI21X1 U1579 ( .A(n5739), .B(n5804), .C(n4003), .Y(n2372) );
  OAI21X1 U1581 ( .A(n5738), .B(n5805), .C(n3913), .Y(n2373) );
  OAI21X1 U1583 ( .A(n5737), .B(n5805), .C(n3277), .Y(n2374) );
  OAI21X1 U1585 ( .A(n5736), .B(n5805), .C(n3201), .Y(n2375) );
  OAI21X1 U1587 ( .A(n5735), .B(n5805), .C(n3125), .Y(n2376) );
  OAI21X1 U1589 ( .A(n5734), .B(n5804), .C(n3049), .Y(n2377) );
  OAI21X1 U1591 ( .A(n5733), .B(n5804), .C(n3830), .Y(n2378) );
  OAI21X1 U1593 ( .A(n5732), .B(n5804), .C(n3747), .Y(n2379) );
  OAI21X1 U1595 ( .A(n5731), .B(n5805), .C(n3665), .Y(n2380) );
  OAI21X1 U1597 ( .A(n5749), .B(n5805), .C(n3276), .Y(n2381) );
  OAI21X1 U1599 ( .A(n5750), .B(n5804), .C(n4270), .Y(n2382) );
  OAI21X1 U1601 ( .A(n5751), .B(n5805), .C(n4179), .Y(n2383) );
  OAI21X1 U1603 ( .A(n5752), .B(n5805), .C(n4092), .Y(n2384) );
  OAI21X1 U1605 ( .A(n5753), .B(n5805), .C(n4002), .Y(n2385) );
  OAI21X1 U1607 ( .A(n5754), .B(n5805), .C(n3912), .Y(n2386) );
  OAI21X1 U1609 ( .A(n5755), .B(n5804), .C(n3200), .Y(n2387) );
  OAI21X1 U1611 ( .A(n5756), .B(n5804), .C(n3124), .Y(n2388) );
  OAI21X1 U1613 ( .A(n5757), .B(n5805), .C(n3048), .Y(n2389) );
  OAI21X1 U1615 ( .A(n5758), .B(n5805), .C(n3829), .Y(n2390) );
  OAI21X1 U1617 ( .A(n5759), .B(n5804), .C(n3746), .Y(n2391) );
  OAI21X1 U1619 ( .A(n5760), .B(n5805), .C(n4178), .Y(n2392) );
  OAI21X1 U1621 ( .A(n5761), .B(n5804), .C(n4091), .Y(n2393) );
  OAI21X1 U1623 ( .A(n5762), .B(n5805), .C(n4001), .Y(n2394) );
  OAI21X1 U1625 ( .A(n5763), .B(n5804), .C(n3047), .Y(n2395) );
  OAI21X1 U1627 ( .A(n5764), .B(n5805), .C(n3586), .Y(n2396) );
  OAI21X1 U1629 ( .A(n5765), .B(n5804), .C(n3508), .Y(n2397) );
  OAI21X1 U1631 ( .A(n5766), .B(n5804), .C(n3429), .Y(n2398) );
  OAI21X1 U1633 ( .A(n5767), .B(n5804), .C(n3351), .Y(n2399) );
  OAI21X1 U1635 ( .A(n5768), .B(n5804), .C(n144), .Y(n2400) );
  OAI21X1 U1637 ( .A(n5769), .B(n5804), .C(n3199), .Y(n2401) );
  OAI21X1 U1639 ( .A(n5770), .B(n5804), .C(n3585), .Y(n2402) );
  OAI21X1 U1641 ( .A(n5771), .B(n5804), .C(n3507), .Y(n2403) );
  OAI21X1 U1643 ( .A(n5772), .B(n5805), .C(n3123), .Y(n2404) );
  OAI21X1 U1645 ( .A(n5748), .B(n5804), .C(n3350), .Y(n2405) );
  OAI21X1 U1647 ( .A(n5747), .B(n5804), .C(n143), .Y(n2406) );
  OAI21X1 U1650 ( .A(n5746), .B(n5802), .C(n3828), .Y(n2407) );
  OAI21X1 U1652 ( .A(n5745), .B(n5802), .C(n3911), .Y(n2408) );
  OAI21X1 U1654 ( .A(n5744), .B(n5802), .C(n3664), .Y(n2409) );
  OAI21X1 U1656 ( .A(n5743), .B(n5802), .C(n3745), .Y(n2410) );
  OAI21X1 U1658 ( .A(n5742), .B(n5803), .C(n4177), .Y(n2411) );
  OAI21X1 U1660 ( .A(n5741), .B(n5802), .C(n4269), .Y(n2412) );
  OAI21X1 U1662 ( .A(n5740), .B(n5803), .C(n4000), .Y(n2413) );
  OAI21X1 U1664 ( .A(n5739), .B(n5802), .C(n4090), .Y(n2414) );
  OAI21X1 U1666 ( .A(n5738), .B(n5803), .C(n3827), .Y(n2415) );
  OAI21X1 U1668 ( .A(n5737), .B(n5803), .C(n3198), .Y(n2416) );
  OAI21X1 U1670 ( .A(n5736), .B(n5803), .C(n3275), .Y(n2417) );
  OAI21X1 U1672 ( .A(n5735), .B(n5803), .C(n3046), .Y(n2418) );
  OAI21X1 U1674 ( .A(n5734), .B(n5802), .C(n3122), .Y(n2419) );
  OAI21X1 U1676 ( .A(n5733), .B(n5802), .C(n3910), .Y(n2420) );
  OAI21X1 U1678 ( .A(n5732), .B(n5802), .C(n3663), .Y(n2421) );
  OAI21X1 U1680 ( .A(n5731), .B(n5803), .C(n3744), .Y(n2422) );
  OAI21X1 U1682 ( .A(n5749), .B(n5803), .C(n3197), .Y(n2423) );
  OAI21X1 U1684 ( .A(n5750), .B(n5802), .C(n4176), .Y(n2424) );
  OAI21X1 U1686 ( .A(n5751), .B(n5803), .C(n4268), .Y(n2425) );
  OAI21X1 U1688 ( .A(n5752), .B(n5803), .C(n3999), .Y(n2426) );
  OAI21X1 U1690 ( .A(n5753), .B(n5803), .C(n4089), .Y(n2427) );
  OAI21X1 U1692 ( .A(n5754), .B(n5803), .C(n3826), .Y(n2428) );
  OAI21X1 U1694 ( .A(n5755), .B(n5802), .C(n3274), .Y(n2429) );
  OAI21X1 U1696 ( .A(n5756), .B(n5802), .C(n3045), .Y(n2430) );
  OAI21X1 U1698 ( .A(n5757), .B(n5803), .C(n3121), .Y(n2431) );
  OAI21X1 U1700 ( .A(n5758), .B(n5803), .C(n3909), .Y(n2432) );
  OAI21X1 U1702 ( .A(n5759), .B(n5802), .C(n3662), .Y(n2433) );
  OAI21X1 U1704 ( .A(n5760), .B(n5803), .C(n4267), .Y(n2434) );
  OAI21X1 U1706 ( .A(n5761), .B(n5802), .C(n3998), .Y(n2435) );
  OAI21X1 U1708 ( .A(n5762), .B(n5803), .C(n4088), .Y(n2436) );
  OAI21X1 U1710 ( .A(n5763), .B(n5802), .C(n3120), .Y(n2437) );
  OAI21X1 U1712 ( .A(n5764), .B(n5803), .C(n3506), .Y(n2438) );
  OAI21X1 U1714 ( .A(n5765), .B(n5802), .C(n3584), .Y(n2439) );
  OAI21X1 U1716 ( .A(n5766), .B(n5802), .C(n3349), .Y(n2440) );
  OAI21X1 U1718 ( .A(n5767), .B(n5802), .C(n3428), .Y(n2441) );
  OAI21X1 U1720 ( .A(n5768), .B(n5802), .C(n142), .Y(n2442) );
  OAI21X1 U1722 ( .A(n5769), .B(n5802), .C(n3273), .Y(n2443) );
  OAI21X1 U1724 ( .A(n5770), .B(n5802), .C(n3505), .Y(n2444) );
  OAI21X1 U1726 ( .A(n5771), .B(n5802), .C(n3583), .Y(n2445) );
  OAI21X1 U1728 ( .A(n5772), .B(n5803), .C(n3044), .Y(n2446) );
  OAI21X1 U1730 ( .A(n5748), .B(n5802), .C(n3427), .Y(n2447) );
  OAI21X1 U1732 ( .A(n5747), .B(n5802), .C(n141), .Y(n2448) );
  OAI21X1 U1735 ( .A(n5746), .B(n5800), .C(n3743), .Y(n2449) );
  OAI21X1 U1737 ( .A(n5745), .B(n5800), .C(n3661), .Y(n2450) );
  OAI21X1 U1739 ( .A(n5744), .B(n5800), .C(n3908), .Y(n2451) );
  OAI21X1 U1741 ( .A(n5743), .B(n5800), .C(n3825), .Y(n2452) );
  OAI21X1 U1743 ( .A(n5742), .B(n5801), .C(n4087), .Y(n2453) );
  OAI21X1 U1745 ( .A(n5741), .B(n5800), .C(n3997), .Y(n2454) );
  OAI21X1 U1747 ( .A(n5740), .B(n5801), .C(n4266), .Y(n2455) );
  OAI21X1 U1749 ( .A(n5739), .B(n5800), .C(n4175), .Y(n2456) );
  OAI21X1 U1751 ( .A(n5738), .B(n5801), .C(n3742), .Y(n2457) );
  OAI21X1 U1753 ( .A(n5737), .B(n5801), .C(n3119), .Y(n2458) );
  OAI21X1 U1755 ( .A(n5736), .B(n5801), .C(n3043), .Y(n2459) );
  OAI21X1 U1757 ( .A(n5735), .B(n5801), .C(n3272), .Y(n2460) );
  OAI21X1 U1759 ( .A(n5734), .B(n5800), .C(n3196), .Y(n2461) );
  OAI21X1 U1761 ( .A(n5733), .B(n5800), .C(n3660), .Y(n2462) );
  OAI21X1 U1763 ( .A(n5732), .B(n5800), .C(n3907), .Y(n2463) );
  OAI21X1 U1765 ( .A(n5731), .B(n5801), .C(n3824), .Y(n2464) );
  OAI21X1 U1767 ( .A(n5749), .B(n5801), .C(n3118), .Y(n2465) );
  OAI21X1 U1769 ( .A(n5750), .B(n5800), .C(n4086), .Y(n2466) );
  OAI21X1 U1771 ( .A(n5751), .B(n5801), .C(n3996), .Y(n2467) );
  OAI21X1 U1773 ( .A(n5752), .B(n5801), .C(n4265), .Y(n2468) );
  OAI21X1 U1775 ( .A(n5753), .B(n5801), .C(n4174), .Y(n2469) );
  OAI21X1 U1777 ( .A(n5754), .B(n5801), .C(n3741), .Y(n2470) );
  OAI21X1 U1779 ( .A(n5755), .B(n5800), .C(n3042), .Y(n2471) );
  OAI21X1 U1781 ( .A(n5756), .B(n5800), .C(n3271), .Y(n2472) );
  OAI21X1 U1783 ( .A(n5757), .B(n5801), .C(n3195), .Y(n2473) );
  OAI21X1 U1785 ( .A(n5758), .B(n5801), .C(n3659), .Y(n2474) );
  OAI21X1 U1787 ( .A(n5759), .B(n5800), .C(n3906), .Y(n2475) );
  OAI21X1 U1789 ( .A(n5760), .B(n5801), .C(n3995), .Y(n2476) );
  OAI21X1 U1791 ( .A(n5761), .B(n5800), .C(n4264), .Y(n2477) );
  OAI21X1 U1793 ( .A(n5762), .B(n5801), .C(n4173), .Y(n2478) );
  OAI21X1 U1795 ( .A(n5763), .B(n5800), .C(n3194), .Y(n2479) );
  OAI21X1 U1797 ( .A(n5764), .B(n5801), .C(n3426), .Y(n2480) );
  OAI21X1 U1799 ( .A(n5765), .B(n5800), .C(n3348), .Y(n2481) );
  OAI21X1 U1801 ( .A(n5766), .B(n5800), .C(n3582), .Y(n2482) );
  OAI21X1 U1803 ( .A(n5767), .B(n5800), .C(n3504), .Y(n2483) );
  OAI21X1 U1805 ( .A(n5768), .B(n5800), .C(n140), .Y(n2484) );
  OAI21X1 U1807 ( .A(n5769), .B(n5800), .C(n3041), .Y(n2485) );
  OAI21X1 U1809 ( .A(n5770), .B(n5800), .C(n3425), .Y(n2486) );
  OAI21X1 U1811 ( .A(n5771), .B(n5800), .C(n3347), .Y(n2487) );
  OAI21X1 U1813 ( .A(n5772), .B(n5801), .C(n3270), .Y(n2488) );
  OAI21X1 U1815 ( .A(n5748), .B(n5800), .C(n3503), .Y(n2489) );
  OAI21X1 U1817 ( .A(n5747), .B(n5800), .C(n139), .Y(n2490) );
  OAI21X1 U1820 ( .A(n5746), .B(n5798), .C(n3658), .Y(n2491) );
  OAI21X1 U1822 ( .A(n5745), .B(n5798), .C(n3740), .Y(n2492) );
  OAI21X1 U1824 ( .A(n5744), .B(n5798), .C(n3823), .Y(n2493) );
  OAI21X1 U1826 ( .A(n5743), .B(n5798), .C(n3905), .Y(n2494) );
  OAI21X1 U1828 ( .A(n5742), .B(n5799), .C(n3994), .Y(n2495) );
  OAI21X1 U1830 ( .A(n5741), .B(n5798), .C(n4085), .Y(n2496) );
  OAI21X1 U1832 ( .A(n5740), .B(n5799), .C(n4172), .Y(n2497) );
  OAI21X1 U1834 ( .A(n5739), .B(n5798), .C(n4263), .Y(n2498) );
  OAI21X1 U1836 ( .A(n5738), .B(n5799), .C(n3657), .Y(n2499) );
  OAI21X1 U1838 ( .A(n5737), .B(n5799), .C(n3040), .Y(n2500) );
  OAI21X1 U1840 ( .A(n5736), .B(n5799), .C(n3117), .Y(n2501) );
  OAI21X1 U1842 ( .A(n5735), .B(n5799), .C(n3193), .Y(n2502) );
  OAI21X1 U1844 ( .A(n5734), .B(n5798), .C(n3269), .Y(n2503) );
  OAI21X1 U1846 ( .A(n5733), .B(n5798), .C(n3739), .Y(n2504) );
  OAI21X1 U1848 ( .A(n5732), .B(n5798), .C(n3822), .Y(n2505) );
  OAI21X1 U1850 ( .A(n5731), .B(n5799), .C(n3904), .Y(n2506) );
  OAI21X1 U1852 ( .A(n5749), .B(n5799), .C(n3039), .Y(n2507) );
  OAI21X1 U1854 ( .A(n5750), .B(n5798), .C(n3993), .Y(n2508) );
  OAI21X1 U1856 ( .A(n5751), .B(n5799), .C(n4084), .Y(n2509) );
  OAI21X1 U1858 ( .A(n5752), .B(n5799), .C(n4171), .Y(n2510) );
  OAI21X1 U1860 ( .A(n5753), .B(n5799), .C(n4262), .Y(n2511) );
  OAI21X1 U1862 ( .A(n5754), .B(n5799), .C(n3656), .Y(n2512) );
  OAI21X1 U1864 ( .A(n5755), .B(n5798), .C(n3116), .Y(n2513) );
  OAI21X1 U1866 ( .A(n5756), .B(n5798), .C(n3192), .Y(n2514) );
  OAI21X1 U1868 ( .A(n5757), .B(n5799), .C(n3268), .Y(n2515) );
  OAI21X1 U1870 ( .A(n5758), .B(n5799), .C(n3738), .Y(n2516) );
  OAI21X1 U1872 ( .A(n5759), .B(n5798), .C(n3821), .Y(n2517) );
  OAI21X1 U1874 ( .A(n5760), .B(n5799), .C(n4083), .Y(n2518) );
  OAI21X1 U1876 ( .A(n5761), .B(n5798), .C(n4170), .Y(n2519) );
  OAI21X1 U1878 ( .A(n5762), .B(n5799), .C(n4261), .Y(n2520) );
  OAI21X1 U1880 ( .A(n5763), .B(n5798), .C(n3267), .Y(n2521) );
  OAI21X1 U1882 ( .A(n5764), .B(n5799), .C(n3346), .Y(n2522) );
  OAI21X1 U1884 ( .A(n5765), .B(n5798), .C(n3424), .Y(n2523) );
  OAI21X1 U1886 ( .A(n5766), .B(n5798), .C(n3502), .Y(n2524) );
  OAI21X1 U1888 ( .A(n5767), .B(n5798), .C(n3581), .Y(n2525) );
  OAI21X1 U1890 ( .A(n5768), .B(n5798), .C(n138), .Y(n2526) );
  OAI21X1 U1892 ( .A(n5769), .B(n5798), .C(n3115), .Y(n2527) );
  OAI21X1 U1894 ( .A(n5770), .B(n5798), .C(n3345), .Y(n2528) );
  OAI21X1 U1896 ( .A(n5771), .B(n5798), .C(n3423), .Y(n2529) );
  OAI21X1 U1898 ( .A(n5772), .B(n5799), .C(n3191), .Y(n2530) );
  OAI21X1 U1900 ( .A(n5748), .B(n5798), .C(n3580), .Y(n2531) );
  OAI21X1 U1902 ( .A(n5747), .B(n5798), .C(n137), .Y(n2532) );
  OAI21X1 U1905 ( .A(n5746), .B(n5796), .C(n3579), .Y(n2533) );
  OAI21X1 U1907 ( .A(n5745), .B(n5796), .C(n3501), .Y(n2534) );
  OAI21X1 U1909 ( .A(n5744), .B(n5796), .C(n3422), .Y(n2535) );
  OAI21X1 U1911 ( .A(n5743), .B(n5796), .C(n3344), .Y(n2536) );
  OAI21X1 U1913 ( .A(n5742), .B(n5797), .C(n3266), .Y(n2537) );
  OAI21X1 U1915 ( .A(n5741), .B(n5796), .C(n3190), .Y(n2538) );
  OAI21X1 U1917 ( .A(n5740), .B(n5797), .C(n3114), .Y(n2539) );
  OAI21X1 U1919 ( .A(n5739), .B(n5796), .C(n3038), .Y(n2540) );
  OAI21X1 U1921 ( .A(n5738), .B(n5797), .C(n3578), .Y(n2541) );
  OAI21X1 U1923 ( .A(n5737), .B(n5797), .C(n4260), .Y(n2542) );
  OAI21X1 U1925 ( .A(n5736), .B(n5797), .C(n4169), .Y(n2543) );
  OAI21X1 U1927 ( .A(n5735), .B(n5797), .C(n4082), .Y(n2544) );
  OAI21X1 U1929 ( .A(n5734), .B(n5796), .C(n3992), .Y(n2545) );
  OAI21X1 U1931 ( .A(n5733), .B(n5796), .C(n3500), .Y(n2546) );
  OAI21X1 U1933 ( .A(n5732), .B(n5796), .C(n3421), .Y(n2547) );
  OAI21X1 U1935 ( .A(n5731), .B(n5797), .C(n3343), .Y(n2548) );
  OAI21X1 U1937 ( .A(n5749), .B(n5797), .C(n4259), .Y(n2549) );
  OAI21X1 U1939 ( .A(n5750), .B(n5796), .C(n3265), .Y(n2550) );
  OAI21X1 U1941 ( .A(n5751), .B(n5797), .C(n3189), .Y(n2551) );
  OAI21X1 U1943 ( .A(n5752), .B(n5797), .C(n3113), .Y(n2552) );
  OAI21X1 U1945 ( .A(n5753), .B(n5797), .C(n3037), .Y(n2553) );
  OAI21X1 U1947 ( .A(n5754), .B(n5797), .C(n3577), .Y(n2554) );
  OAI21X1 U1949 ( .A(n5755), .B(n5796), .C(n4168), .Y(n2555) );
  OAI21X1 U1951 ( .A(n5756), .B(n5796), .C(n4081), .Y(n2556) );
  OAI21X1 U1953 ( .A(n5757), .B(n5797), .C(n3991), .Y(n2557) );
  OAI21X1 U1955 ( .A(n5758), .B(n5797), .C(n3499), .Y(n2558) );
  OAI21X1 U1957 ( .A(n5759), .B(n5796), .C(n3420), .Y(n2559) );
  OAI21X1 U1959 ( .A(n5760), .B(n5797), .C(n3188), .Y(n2560) );
  OAI21X1 U1961 ( .A(n5761), .B(n5796), .C(n3112), .Y(n2561) );
  OAI21X1 U1963 ( .A(n5762), .B(n5797), .C(n3036), .Y(n2562) );
  OAI21X1 U1965 ( .A(n5763), .B(n5796), .C(n3990), .Y(n2563) );
  OAI21X1 U1967 ( .A(n5764), .B(n5797), .C(n3903), .Y(n2564) );
  OAI21X1 U1969 ( .A(n5765), .B(n5796), .C(n3820), .Y(n2565) );
  OAI21X1 U1971 ( .A(n5766), .B(n5796), .C(n3737), .Y(n2566) );
  OAI21X1 U1973 ( .A(n5767), .B(n5796), .C(n3655), .Y(n2567) );
  OAI21X1 U1975 ( .A(n5768), .B(n5796), .C(n136), .Y(n2568) );
  OAI21X1 U1977 ( .A(n5769), .B(n5796), .C(n4167), .Y(n2569) );
  OAI21X1 U1979 ( .A(n5770), .B(n5796), .C(n3902), .Y(n2570) );
  OAI21X1 U1981 ( .A(n5771), .B(n5796), .C(n3819), .Y(n2571) );
  OAI21X1 U1983 ( .A(n5772), .B(n5797), .C(n4080), .Y(n2572) );
  OAI21X1 U1985 ( .A(n5748), .B(n5796), .C(n3654), .Y(n2573) );
  OAI21X1 U1987 ( .A(n5747), .B(n5796), .C(n135), .Y(n2574) );
  OAI21X1 U1990 ( .A(n5746), .B(n5794), .C(n3498), .Y(n2575) );
  OAI21X1 U1992 ( .A(n5745), .B(n5794), .C(n3576), .Y(n2576) );
  OAI21X1 U1994 ( .A(n5744), .B(n5794), .C(n3342), .Y(n2577) );
  OAI21X1 U1996 ( .A(n5743), .B(n5794), .C(n3419), .Y(n2578) );
  OAI21X1 U1998 ( .A(n5742), .B(n5795), .C(n3187), .Y(n2579) );
  OAI21X1 U2000 ( .A(n5741), .B(n5794), .C(n3264), .Y(n2580) );
  OAI21X1 U2002 ( .A(n5740), .B(n5795), .C(n3035), .Y(n2581) );
  OAI21X1 U2004 ( .A(n5739), .B(n5794), .C(n3111), .Y(n2582) );
  OAI21X1 U2006 ( .A(n5738), .B(n5795), .C(n3497), .Y(n2583) );
  OAI21X1 U2008 ( .A(n5737), .B(n5795), .C(n4166), .Y(n2584) );
  OAI21X1 U2010 ( .A(n5736), .B(n5795), .C(n4258), .Y(n2585) );
  OAI21X1 U2012 ( .A(n5735), .B(n5795), .C(n3989), .Y(n2586) );
  OAI21X1 U2014 ( .A(n5734), .B(n5794), .C(n4079), .Y(n2587) );
  OAI21X1 U2016 ( .A(n5733), .B(n5794), .C(n3575), .Y(n2588) );
  OAI21X1 U2018 ( .A(n5732), .B(n5794), .C(n3341), .Y(n2589) );
  OAI21X1 U2020 ( .A(n5731), .B(n5795), .C(n3418), .Y(n2590) );
  OAI21X1 U2022 ( .A(n5749), .B(n5795), .C(n4165), .Y(n2591) );
  OAI21X1 U2024 ( .A(n5750), .B(n5794), .C(n3186), .Y(n2592) );
  OAI21X1 U2026 ( .A(n5751), .B(n5795), .C(n3263), .Y(n2593) );
  OAI21X1 U2028 ( .A(n5752), .B(n5795), .C(n3034), .Y(n2594) );
  OAI21X1 U2030 ( .A(n5753), .B(n5795), .C(n3110), .Y(n2595) );
  OAI21X1 U2032 ( .A(n5754), .B(n5795), .C(n3496), .Y(n2596) );
  OAI21X1 U2034 ( .A(n5755), .B(n5794), .C(n4257), .Y(n2597) );
  OAI21X1 U2036 ( .A(n5756), .B(n5794), .C(n3988), .Y(n2598) );
  OAI21X1 U2038 ( .A(n5757), .B(n5795), .C(n4078), .Y(n2599) );
  OAI21X1 U2040 ( .A(n5758), .B(n5795), .C(n3574), .Y(n2600) );
  OAI21X1 U2042 ( .A(n5759), .B(n5794), .C(n3340), .Y(n2601) );
  OAI21X1 U2044 ( .A(n5760), .B(n5795), .C(n3262), .Y(n2602) );
  OAI21X1 U2046 ( .A(n5761), .B(n5794), .C(n3033), .Y(n2603) );
  OAI21X1 U2048 ( .A(n5762), .B(n5795), .C(n3109), .Y(n2604) );
  OAI21X1 U2050 ( .A(n5763), .B(n5794), .C(n4077), .Y(n2605) );
  OAI21X1 U2052 ( .A(n5764), .B(n5795), .C(n3818), .Y(n2606) );
  OAI21X1 U2054 ( .A(n5765), .B(n5794), .C(n3901), .Y(n2607) );
  OAI21X1 U2056 ( .A(n5766), .B(n5794), .C(n3653), .Y(n2608) );
  OAI21X1 U2058 ( .A(n5767), .B(n5794), .C(n3736), .Y(n2609) );
  OAI21X1 U2060 ( .A(n5768), .B(n5794), .C(n134), .Y(n2610) );
  OAI21X1 U2062 ( .A(n5769), .B(n5794), .C(n4256), .Y(n2611) );
  OAI21X1 U2064 ( .A(n5770), .B(n5794), .C(n3817), .Y(n2612) );
  OAI21X1 U2066 ( .A(n5771), .B(n5794), .C(n3900), .Y(n2613) );
  OAI21X1 U2068 ( .A(n5772), .B(n5795), .C(n3987), .Y(n2614) );
  OAI21X1 U2070 ( .A(n5748), .B(n5794), .C(n3735), .Y(n2615) );
  OAI21X1 U2072 ( .A(n5747), .B(n5794), .C(n133), .Y(n2616) );
  OAI21X1 U2075 ( .A(n5746), .B(n5792), .C(n3417), .Y(n2617) );
  OAI21X1 U2077 ( .A(n5745), .B(n5792), .C(n3339), .Y(n2618) );
  OAI21X1 U2079 ( .A(n5744), .B(n5792), .C(n3573), .Y(n2619) );
  OAI21X1 U2081 ( .A(n5743), .B(n5792), .C(n3495), .Y(n2620) );
  OAI21X1 U2083 ( .A(n5742), .B(n5793), .C(n3108), .Y(n2621) );
  OAI21X1 U2085 ( .A(n5741), .B(n5792), .C(n3032), .Y(n2622) );
  OAI21X1 U2087 ( .A(n5740), .B(n5793), .C(n3261), .Y(n2623) );
  OAI21X1 U2089 ( .A(n5739), .B(n5792), .C(n3185), .Y(n2624) );
  OAI21X1 U2091 ( .A(n5738), .B(n5793), .C(n3416), .Y(n2625) );
  OAI21X1 U2093 ( .A(n5737), .B(n5793), .C(n4076), .Y(n2626) );
  OAI21X1 U2095 ( .A(n5736), .B(n5793), .C(n3986), .Y(n2627) );
  OAI21X1 U2097 ( .A(n5735), .B(n5793), .C(n4255), .Y(n2628) );
  OAI21X1 U2099 ( .A(n5734), .B(n5792), .C(n4164), .Y(n2629) );
  OAI21X1 U2101 ( .A(n5733), .B(n5792), .C(n3338), .Y(n2630) );
  OAI21X1 U2103 ( .A(n5732), .B(n5792), .C(n3572), .Y(n2631) );
  OAI21X1 U2105 ( .A(n5731), .B(n5793), .C(n3494), .Y(n2632) );
  OAI21X1 U2107 ( .A(n5749), .B(n5793), .C(n4075), .Y(n2633) );
  OAI21X1 U2109 ( .A(n5750), .B(n5792), .C(n3107), .Y(n2634) );
  OAI21X1 U2111 ( .A(n5751), .B(n5793), .C(n3031), .Y(n2635) );
  OAI21X1 U2113 ( .A(n5752), .B(n5793), .C(n3260), .Y(n2636) );
  OAI21X1 U2115 ( .A(n5753), .B(n5793), .C(n3184), .Y(n2637) );
  OAI21X1 U2117 ( .A(n5754), .B(n5793), .C(n3415), .Y(n2638) );
  OAI21X1 U2119 ( .A(n5755), .B(n5792), .C(n3985), .Y(n2639) );
  OAI21X1 U2121 ( .A(n5756), .B(n5792), .C(n4254), .Y(n2640) );
  OAI21X1 U2123 ( .A(n5757), .B(n5793), .C(n4163), .Y(n2641) );
  OAI21X1 U2125 ( .A(n5758), .B(n5793), .C(n3337), .Y(n2642) );
  OAI21X1 U2127 ( .A(n5759), .B(n5792), .C(n3571), .Y(n2643) );
  OAI21X1 U2129 ( .A(n5760), .B(n5793), .C(n3030), .Y(n2644) );
  OAI21X1 U2131 ( .A(n5761), .B(n5792), .C(n3259), .Y(n2645) );
  OAI21X1 U2133 ( .A(n5762), .B(n5793), .C(n3183), .Y(n2646) );
  OAI21X1 U2135 ( .A(n5763), .B(n5792), .C(n4162), .Y(n2647) );
  OAI21X1 U2137 ( .A(n5764), .B(n5793), .C(n3734), .Y(n2648) );
  OAI21X1 U2139 ( .A(n5765), .B(n5792), .C(n3652), .Y(n2649) );
  OAI21X1 U2141 ( .A(n5766), .B(n5792), .C(n3899), .Y(n2650) );
  OAI21X1 U2143 ( .A(n5767), .B(n5792), .C(n3816), .Y(n2651) );
  OAI21X1 U2145 ( .A(n5768), .B(n5792), .C(n132), .Y(n2652) );
  OAI21X1 U2147 ( .A(n5769), .B(n5792), .C(n3984), .Y(n2653) );
  OAI21X1 U2149 ( .A(n5770), .B(n5792), .C(n3733), .Y(n2654) );
  OAI21X1 U2151 ( .A(n5771), .B(n5792), .C(n3651), .Y(n2655) );
  OAI21X1 U2153 ( .A(n5772), .B(n5793), .C(n4253), .Y(n2656) );
  OAI21X1 U2155 ( .A(n5748), .B(n5792), .C(n3815), .Y(n2657) );
  OAI21X1 U2157 ( .A(n5747), .B(n5792), .C(n131), .Y(n2658) );
  NOR3X1 U2160 ( .A(n1568), .B(wr_ptr[3]), .C(n5902), .Y(n919) );
  OAI21X1 U2161 ( .A(n5746), .B(n5791), .C(n3336), .Y(n2659) );
  OAI21X1 U2163 ( .A(n5745), .B(n5790), .C(n3414), .Y(n2660) );
  OAI21X1 U2165 ( .A(n5744), .B(n5790), .C(n3493), .Y(n2661) );
  OAI21X1 U2167 ( .A(n5743), .B(n5790), .C(n3570), .Y(n2662) );
  OAI21X1 U2169 ( .A(n5742), .B(n5790), .C(n3029), .Y(n2663) );
  OAI21X1 U2171 ( .A(n5741), .B(n5790), .C(n3106), .Y(n2664) );
  OAI21X1 U2173 ( .A(n5740), .B(n5790), .C(n3182), .Y(n2665) );
  OAI21X1 U2175 ( .A(n5739), .B(n5790), .C(n3258), .Y(n2666) );
  OAI21X1 U2177 ( .A(n5738), .B(n5790), .C(n3335), .Y(n2667) );
  OAI21X1 U2179 ( .A(n5737), .B(n5790), .C(n3983), .Y(n2668) );
  OAI21X1 U2181 ( .A(n5736), .B(n5790), .C(n4074), .Y(n2669) );
  OAI21X1 U2183 ( .A(n5735), .B(n5790), .C(n4161), .Y(n2670) );
  OAI21X1 U2185 ( .A(n5734), .B(n5790), .C(n4252), .Y(n2671) );
  OAI21X1 U2187 ( .A(n5733), .B(n5790), .C(n3413), .Y(n2672) );
  OAI21X1 U2189 ( .A(n5732), .B(n5790), .C(n3492), .Y(n2673) );
  OAI21X1 U2191 ( .A(n5731), .B(n5791), .C(n3569), .Y(n2674) );
  OAI21X1 U2193 ( .A(n5749), .B(n5791), .C(n3982), .Y(n2675) );
  OAI21X1 U2195 ( .A(n5750), .B(n5790), .C(n3028), .Y(n2676) );
  OAI21X1 U2197 ( .A(n5751), .B(n5791), .C(n3105), .Y(n2677) );
  OAI21X1 U2199 ( .A(n5752), .B(n5790), .C(n3181), .Y(n2678) );
  OAI21X1 U2201 ( .A(n5753), .B(n5790), .C(n3257), .Y(n2679) );
  OAI21X1 U2203 ( .A(n5754), .B(n5791), .C(n3334), .Y(n2680) );
  OAI21X1 U2205 ( .A(n5755), .B(n5790), .C(n4073), .Y(n2681) );
  OAI21X1 U2207 ( .A(n5756), .B(n5790), .C(n4160), .Y(n2682) );
  OAI21X1 U2209 ( .A(n5757), .B(n5790), .C(n4251), .Y(n2683) );
  OAI21X1 U2211 ( .A(n5758), .B(n5791), .C(n3412), .Y(n2684) );
  OAI21X1 U2213 ( .A(n5759), .B(n5790), .C(n3491), .Y(n2685) );
  OAI21X1 U2215 ( .A(n5760), .B(n5790), .C(n3104), .Y(n2686) );
  OAI21X1 U2217 ( .A(n5761), .B(n5791), .C(n3180), .Y(n2687) );
  OAI21X1 U2219 ( .A(n5762), .B(n5791), .C(n3256), .Y(n2688) );
  OAI21X1 U2221 ( .A(n5763), .B(n5790), .C(n4250), .Y(n2689) );
  OAI21X1 U2223 ( .A(n5764), .B(n5790), .C(n3650), .Y(n2690) );
  OAI21X1 U2225 ( .A(n5765), .B(n5791), .C(n3732), .Y(n2691) );
  OAI21X1 U2227 ( .A(n5766), .B(n5791), .C(n3814), .Y(n2692) );
  OAI21X1 U2229 ( .A(n5767), .B(n5790), .C(n3898), .Y(n2693) );
  OAI21X1 U2231 ( .A(n5768), .B(n5791), .C(n130), .Y(n2694) );
  OAI21X1 U2233 ( .A(n5769), .B(n5790), .C(n4072), .Y(n2695) );
  OAI21X1 U2235 ( .A(n5770), .B(n5790), .C(n3649), .Y(n2696) );
  OAI21X1 U2237 ( .A(n5771), .B(n5791), .C(n3731), .Y(n2697) );
  OAI21X1 U2239 ( .A(n5772), .B(n5791), .C(n4159), .Y(n2698) );
  OAI21X1 U2241 ( .A(n5748), .B(n5791), .C(n3897), .Y(n2699) );
  OAI21X1 U2243 ( .A(n5747), .B(n5790), .C(n129), .Y(n2700) );
  NOR3X1 U2246 ( .A(wr_ptr[1]), .B(wr_ptr[2]), .C(wr_ptr[0]), .Y(n221) );
  OAI21X1 U2247 ( .A(n5746), .B(n5789), .C(n3255), .Y(n2701) );
  OAI21X1 U2249 ( .A(n5745), .B(n5788), .C(n3179), .Y(n2702) );
  OAI21X1 U2251 ( .A(n5744), .B(n5788), .C(n3103), .Y(n2703) );
  OAI21X1 U2253 ( .A(n5743), .B(n5788), .C(n3027), .Y(n2704) );
  OAI21X1 U2255 ( .A(n5742), .B(n5788), .C(n3568), .Y(n2705) );
  OAI21X1 U2257 ( .A(n5741), .B(n5788), .C(n3490), .Y(n2706) );
  OAI21X1 U2259 ( .A(n5740), .B(n5788), .C(n3411), .Y(n2707) );
  OAI21X1 U2261 ( .A(n5739), .B(n5788), .C(n3333), .Y(n2708) );
  OAI21X1 U2263 ( .A(n5738), .B(n5788), .C(n3254), .Y(n2709) );
  OAI21X1 U2265 ( .A(n5737), .B(n5788), .C(n3896), .Y(n2710) );
  OAI21X1 U2267 ( .A(n5736), .B(n5788), .C(n3813), .Y(n2711) );
  OAI21X1 U2269 ( .A(n5735), .B(n5788), .C(n3730), .Y(n2712) );
  OAI21X1 U2271 ( .A(n5734), .B(n5788), .C(n3648), .Y(n2713) );
  OAI21X1 U2273 ( .A(n5733), .B(n5788), .C(n3178), .Y(n2714) );
  OAI21X1 U2275 ( .A(n5732), .B(n5788), .C(n3102), .Y(n2715) );
  OAI21X1 U2277 ( .A(n5731), .B(n5789), .C(n3026), .Y(n2716) );
  OAI21X1 U2279 ( .A(n5749), .B(n5789), .C(n3895), .Y(n2717) );
  OAI21X1 U2281 ( .A(n5750), .B(n5788), .C(n3567), .Y(n2718) );
  OAI21X1 U2283 ( .A(n5751), .B(n5789), .C(n3489), .Y(n2719) );
  OAI21X1 U2285 ( .A(n5752), .B(n5788), .C(n3410), .Y(n2720) );
  OAI21X1 U2287 ( .A(n5753), .B(n5788), .C(n3332), .Y(n2721) );
  OAI21X1 U2289 ( .A(n5754), .B(n5789), .C(n3253), .Y(n2722) );
  OAI21X1 U2291 ( .A(n5755), .B(n5788), .C(n3812), .Y(n2723) );
  OAI21X1 U2293 ( .A(n5756), .B(n5788), .C(n3729), .Y(n2724) );
  OAI21X1 U2295 ( .A(n5757), .B(n5788), .C(n3647), .Y(n2725) );
  OAI21X1 U2297 ( .A(n5758), .B(n5789), .C(n3177), .Y(n2726) );
  OAI21X1 U2299 ( .A(n5759), .B(n5788), .C(n3101), .Y(n2727) );
  OAI21X1 U2301 ( .A(n5760), .B(n5788), .C(n3488), .Y(n2728) );
  OAI21X1 U2303 ( .A(n5761), .B(n5789), .C(n3409), .Y(n2729) );
  OAI21X1 U2305 ( .A(n5762), .B(n5789), .C(n3331), .Y(n2730) );
  OAI21X1 U2307 ( .A(n5763), .B(n5788), .C(n3646), .Y(n2731) );
  OAI21X1 U2309 ( .A(n5764), .B(n5788), .C(n4249), .Y(n2732) );
  OAI21X1 U2311 ( .A(n5765), .B(n5789), .C(n4158), .Y(n2733) );
  OAI21X1 U2313 ( .A(n5766), .B(n5789), .C(n4071), .Y(n2734) );
  OAI21X1 U2315 ( .A(n5767), .B(n5788), .C(n3981), .Y(n2735) );
  OAI21X1 U2317 ( .A(n5768), .B(n5789), .C(n128), .Y(n2736) );
  OAI21X1 U2319 ( .A(n5769), .B(n5788), .C(n3811), .Y(n2737) );
  OAI21X1 U2321 ( .A(n5770), .B(n5788), .C(n4248), .Y(n2738) );
  OAI21X1 U2323 ( .A(n5771), .B(n5789), .C(n4157), .Y(n2739) );
  OAI21X1 U2325 ( .A(n5772), .B(n5789), .C(n3728), .Y(n2740) );
  OAI21X1 U2327 ( .A(n5748), .B(n5789), .C(n3980), .Y(n2741) );
  OAI21X1 U2329 ( .A(n5747), .B(n5788), .C(n127), .Y(n2742) );
  NOR3X1 U2332 ( .A(wr_ptr[1]), .B(wr_ptr[2]), .C(n5898), .Y(n266) );
  OAI21X1 U2333 ( .A(n5746), .B(n5786), .C(n4247), .Y(n2743) );
  OAI21X1 U2335 ( .A(n5745), .B(n5786), .C(n4156), .Y(n2744) );
  OAI21X1 U2337 ( .A(n5744), .B(n5786), .C(n4070), .Y(n2745) );
  OAI21X1 U2339 ( .A(n5743), .B(n5787), .C(n3979), .Y(n2746) );
  OAI21X1 U2341 ( .A(n5742), .B(n5786), .C(n3894), .Y(n2747) );
  OAI21X1 U2343 ( .A(n5741), .B(n5787), .C(n3810), .Y(n2748) );
  OAI21X1 U2345 ( .A(n5740), .B(n5787), .C(n3727), .Y(n2749) );
  OAI21X1 U2347 ( .A(n5739), .B(n5787), .C(n3645), .Y(n2750) );
  OAI21X1 U2349 ( .A(n5738), .B(n5786), .C(n4246), .Y(n2751) );
  OAI21X1 U2351 ( .A(n5737), .B(n5786), .C(n3566), .Y(n2752) );
  OAI21X1 U2353 ( .A(n5736), .B(n5787), .C(n3487), .Y(n2753) );
  OAI21X1 U2355 ( .A(n5735), .B(n5786), .C(n3408), .Y(n2754) );
  OAI21X1 U2357 ( .A(n5734), .B(n5787), .C(n3330), .Y(n2755) );
  OAI21X1 U2359 ( .A(n5733), .B(n5786), .C(n4155), .Y(n2756) );
  OAI21X1 U2361 ( .A(n5732), .B(n5787), .C(n4069), .Y(n2757) );
  OAI21X1 U2363 ( .A(n5731), .B(n5786), .C(n3978), .Y(n2758) );
  OAI21X1 U2365 ( .A(n5749), .B(n5787), .C(n3565), .Y(n2759) );
  OAI21X1 U2367 ( .A(n5750), .B(n5786), .C(n3893), .Y(n2760) );
  OAI21X1 U2369 ( .A(n5751), .B(n5786), .C(n3809), .Y(n2761) );
  OAI21X1 U2371 ( .A(n5752), .B(n5787), .C(n3726), .Y(n2762) );
  OAI21X1 U2373 ( .A(n5753), .B(n5786), .C(n3644), .Y(n2763) );
  OAI21X1 U2375 ( .A(n5754), .B(n5786), .C(n4245), .Y(n2764) );
  OAI21X1 U2377 ( .A(n5755), .B(n5787), .C(n3486), .Y(n2765) );
  OAI21X1 U2379 ( .A(n5756), .B(n5787), .C(n3407), .Y(n2766) );
  OAI21X1 U2381 ( .A(n5757), .B(n5786), .C(n3329), .Y(n2767) );
  OAI21X1 U2383 ( .A(n5758), .B(n5787), .C(n4154), .Y(n2768) );
  OAI21X1 U2385 ( .A(n5759), .B(n5786), .C(n4068), .Y(n2769) );
  OAI21X1 U2387 ( .A(n5760), .B(n5786), .C(n3808), .Y(n2770) );
  OAI21X1 U2389 ( .A(n5761), .B(n5787), .C(n3725), .Y(n2771) );
  OAI21X1 U2391 ( .A(n5762), .B(n5787), .C(n3643), .Y(n2772) );
  OAI21X1 U2393 ( .A(n5763), .B(n5787), .C(n3328), .Y(n2773) );
  OAI21X1 U2395 ( .A(n5764), .B(n5786), .C(n3252), .Y(n2774) );
  OAI21X1 U2397 ( .A(n5765), .B(n5787), .C(n3176), .Y(n2775) );
  OAI21X1 U2399 ( .A(n5766), .B(n5787), .C(n3100), .Y(n2776) );
  OAI21X1 U2401 ( .A(n5767), .B(n5787), .C(n3025), .Y(n2777) );
  OAI21X1 U2403 ( .A(n5768), .B(n5786), .C(n126), .Y(n2778) );
  OAI21X1 U2405 ( .A(n5769), .B(n5787), .C(n3485), .Y(n2779) );
  OAI21X1 U2407 ( .A(n5770), .B(n5786), .C(n3251), .Y(n2780) );
  OAI21X1 U2409 ( .A(n5771), .B(n5787), .C(n3175), .Y(n2781) );
  OAI21X1 U2411 ( .A(n5772), .B(n5786), .C(n3406), .Y(n2782) );
  OAI21X1 U2413 ( .A(n5748), .B(n5787), .C(n3024), .Y(n2783) );
  OAI21X1 U2415 ( .A(n5747), .B(n5786), .C(n125), .Y(n2784) );
  NOR3X1 U2418 ( .A(wr_ptr[0]), .B(wr_ptr[2]), .C(n5899), .Y(n310) );
  OAI21X1 U2419 ( .A(n5746), .B(n5784), .C(n4153), .Y(n2785) );
  OAI21X1 U2421 ( .A(n5745), .B(n5784), .C(n4244), .Y(n2786) );
  OAI21X1 U2423 ( .A(n5744), .B(n5784), .C(n3977), .Y(n2787) );
  OAI21X1 U2425 ( .A(n5743), .B(n5785), .C(n4067), .Y(n2788) );
  OAI21X1 U2427 ( .A(n5742), .B(n5784), .C(n3807), .Y(n2789) );
  OAI21X1 U2429 ( .A(n5741), .B(n5785), .C(n3892), .Y(n2790) );
  OAI21X1 U2431 ( .A(n5740), .B(n5785), .C(n3642), .Y(n2791) );
  OAI21X1 U2433 ( .A(n5739), .B(n5785), .C(n3724), .Y(n2792) );
  OAI21X1 U2435 ( .A(n5738), .B(n5784), .C(n4152), .Y(n2793) );
  OAI21X1 U2437 ( .A(n5737), .B(n5784), .C(n3484), .Y(n2794) );
  OAI21X1 U2439 ( .A(n5736), .B(n5785), .C(n3564), .Y(n2795) );
  OAI21X1 U2441 ( .A(n5735), .B(n5784), .C(n3327), .Y(n2796) );
  OAI21X1 U2443 ( .A(n5734), .B(n5785), .C(n3405), .Y(n2797) );
  OAI21X1 U2445 ( .A(n5733), .B(n5784), .C(n4243), .Y(n2798) );
  OAI21X1 U2447 ( .A(n5732), .B(n5785), .C(n3976), .Y(n2799) );
  OAI21X1 U2449 ( .A(n5731), .B(n5784), .C(n4066), .Y(n2800) );
  OAI21X1 U2451 ( .A(n5749), .B(n5785), .C(n3483), .Y(n2801) );
  OAI21X1 U2453 ( .A(n5750), .B(n5784), .C(n3806), .Y(n2802) );
  OAI21X1 U2455 ( .A(n5751), .B(n5784), .C(n3891), .Y(n2803) );
  OAI21X1 U2457 ( .A(n5752), .B(n5785), .C(n3641), .Y(n2804) );
  OAI21X1 U2459 ( .A(n5753), .B(n5784), .C(n3723), .Y(n2805) );
  OAI21X1 U2461 ( .A(n5754), .B(n5784), .C(n4151), .Y(n2806) );
  OAI21X1 U2463 ( .A(n5755), .B(n5785), .C(n3563), .Y(n2807) );
  OAI21X1 U2465 ( .A(n5756), .B(n5785), .C(n3326), .Y(n2808) );
  OAI21X1 U2467 ( .A(n5757), .B(n5784), .C(n3404), .Y(n2809) );
  OAI21X1 U2469 ( .A(n5758), .B(n5785), .C(n4242), .Y(n2810) );
  OAI21X1 U2471 ( .A(n5759), .B(n5784), .C(n3975), .Y(n2811) );
  OAI21X1 U2473 ( .A(n5760), .B(n5784), .C(n3890), .Y(n2812) );
  OAI21X1 U2475 ( .A(n5761), .B(n5785), .C(n3640), .Y(n2813) );
  OAI21X1 U2477 ( .A(n5762), .B(n5785), .C(n3722), .Y(n2814) );
  OAI21X1 U2479 ( .A(n5763), .B(n5785), .C(n3403), .Y(n2815) );
  OAI21X1 U2481 ( .A(n5764), .B(n5784), .C(n3174), .Y(n2816) );
  OAI21X1 U2483 ( .A(n5765), .B(n5785), .C(n3250), .Y(n2817) );
  OAI21X1 U2485 ( .A(n5766), .B(n5785), .C(n3023), .Y(n2818) );
  OAI21X1 U2487 ( .A(n5767), .B(n5785), .C(n3099), .Y(n2819) );
  OAI21X1 U2489 ( .A(n5768), .B(n5784), .C(n124), .Y(n2820) );
  OAI21X1 U2491 ( .A(n5769), .B(n5785), .C(n3562), .Y(n2821) );
  OAI21X1 U2493 ( .A(n5770), .B(n5784), .C(n3173), .Y(n2822) );
  OAI21X1 U2495 ( .A(n5771), .B(n5785), .C(n3249), .Y(n2823) );
  OAI21X1 U2497 ( .A(n5772), .B(n5784), .C(n3325), .Y(n2824) );
  OAI21X1 U2499 ( .A(n5748), .B(n5785), .C(n3098), .Y(n2825) );
  OAI21X1 U2501 ( .A(n5747), .B(n5784), .C(n123), .Y(n2826) );
  NOR3X1 U2504 ( .A(n5898), .B(wr_ptr[2]), .C(n5899), .Y(n354) );
  OAI21X1 U2505 ( .A(n5746), .B(n5782), .C(n4065), .Y(n2827) );
  OAI21X1 U2507 ( .A(n5745), .B(n5782), .C(n3974), .Y(n2828) );
  OAI21X1 U2509 ( .A(n5744), .B(n5782), .C(n4241), .Y(n2829) );
  OAI21X1 U2511 ( .A(n5743), .B(n5783), .C(n4150), .Y(n2830) );
  OAI21X1 U2513 ( .A(n5742), .B(n5782), .C(n3721), .Y(n2831) );
  OAI21X1 U2515 ( .A(n5741), .B(n5783), .C(n3639), .Y(n2832) );
  OAI21X1 U2517 ( .A(n5740), .B(n5783), .C(n3889), .Y(n2833) );
  OAI21X1 U2519 ( .A(n5739), .B(n5783), .C(n3805), .Y(n2834) );
  OAI21X1 U2521 ( .A(n5738), .B(n5782), .C(n4064), .Y(n2835) );
  OAI21X1 U2523 ( .A(n5737), .B(n5782), .C(n3402), .Y(n2836) );
  OAI21X1 U2525 ( .A(n5736), .B(n5783), .C(n3324), .Y(n2837) );
  OAI21X1 U2527 ( .A(n5735), .B(n5782), .C(n3561), .Y(n2838) );
  OAI21X1 U2529 ( .A(n5734), .B(n5783), .C(n3482), .Y(n2839) );
  OAI21X1 U2531 ( .A(n5733), .B(n5782), .C(n3973), .Y(n2840) );
  OAI21X1 U2533 ( .A(n5732), .B(n5783), .C(n4240), .Y(n2841) );
  OAI21X1 U2535 ( .A(n5731), .B(n5782), .C(n4149), .Y(n2842) );
  OAI21X1 U2537 ( .A(n5749), .B(n5783), .C(n3401), .Y(n2843) );
  OAI21X1 U2539 ( .A(n5750), .B(n5782), .C(n3720), .Y(n2844) );
  OAI21X1 U2541 ( .A(n5751), .B(n5782), .C(n3638), .Y(n2845) );
  OAI21X1 U2543 ( .A(n5752), .B(n5783), .C(n3888), .Y(n2846) );
  OAI21X1 U2545 ( .A(n5753), .B(n5782), .C(n3804), .Y(n2847) );
  OAI21X1 U2547 ( .A(n5754), .B(n5782), .C(n4063), .Y(n2848) );
  OAI21X1 U2549 ( .A(n5755), .B(n5783), .C(n3323), .Y(n2849) );
  OAI21X1 U2551 ( .A(n5756), .B(n5783), .C(n3560), .Y(n2850) );
  OAI21X1 U2553 ( .A(n5757), .B(n5782), .C(n3481), .Y(n2851) );
  OAI21X1 U2555 ( .A(n5758), .B(n5783), .C(n3972), .Y(n2852) );
  OAI21X1 U2557 ( .A(n5759), .B(n5782), .C(n4239), .Y(n2853) );
  OAI21X1 U2559 ( .A(n5760), .B(n5782), .C(n3637), .Y(n2854) );
  OAI21X1 U2561 ( .A(n5761), .B(n5783), .C(n3887), .Y(n2855) );
  OAI21X1 U2563 ( .A(n5762), .B(n5783), .C(n3803), .Y(n2856) );
  OAI21X1 U2565 ( .A(n5763), .B(n5783), .C(n3480), .Y(n2857) );
  OAI21X1 U2567 ( .A(n5764), .B(n5782), .C(n3097), .Y(n2858) );
  OAI21X1 U2569 ( .A(n5765), .B(n5783), .C(n3022), .Y(n2859) );
  OAI21X1 U2571 ( .A(n5766), .B(n5783), .C(n3248), .Y(n2860) );
  OAI21X1 U2573 ( .A(n5767), .B(n5783), .C(n3172), .Y(n2861) );
  OAI21X1 U2575 ( .A(n5768), .B(n5782), .C(n122), .Y(n2862) );
  OAI21X1 U2577 ( .A(n5769), .B(n5783), .C(n3322), .Y(n2863) );
  OAI21X1 U2579 ( .A(n5770), .B(n5782), .C(n3096), .Y(n2864) );
  OAI21X1 U2581 ( .A(n5771), .B(n5783), .C(n3021), .Y(n2865) );
  OAI21X1 U2583 ( .A(n5772), .B(n5782), .C(n3559), .Y(n2866) );
  OAI21X1 U2585 ( .A(n5748), .B(n5783), .C(n3171), .Y(n2867) );
  OAI21X1 U2587 ( .A(n5747), .B(n5782), .C(n121), .Y(n2868) );
  NOR3X1 U2590 ( .A(wr_ptr[0]), .B(wr_ptr[1]), .C(n5900), .Y(n398) );
  OAI21X1 U2591 ( .A(n5746), .B(n5780), .C(n3971), .Y(n2869) );
  OAI21X1 U2593 ( .A(n5745), .B(n5780), .C(n4062), .Y(n2870) );
  OAI21X1 U2595 ( .A(n5744), .B(n5780), .C(n4148), .Y(n2871) );
  OAI21X1 U2597 ( .A(n5743), .B(n5781), .C(n4238), .Y(n2872) );
  OAI21X1 U2599 ( .A(n5742), .B(n5780), .C(n3636), .Y(n2873) );
  OAI21X1 U2601 ( .A(n5741), .B(n5781), .C(n3719), .Y(n2874) );
  OAI21X1 U2603 ( .A(n5740), .B(n5781), .C(n3802), .Y(n2875) );
  OAI21X1 U2605 ( .A(n5739), .B(n5781), .C(n3886), .Y(n2876) );
  OAI21X1 U2607 ( .A(n5738), .B(n5780), .C(n3970), .Y(n2877) );
  OAI21X1 U2609 ( .A(n5737), .B(n5780), .C(n3321), .Y(n2878) );
  OAI21X1 U2611 ( .A(n5736), .B(n5781), .C(n3400), .Y(n2879) );
  OAI21X1 U2613 ( .A(n5735), .B(n5780), .C(n3479), .Y(n2880) );
  OAI21X1 U2615 ( .A(n5734), .B(n5781), .C(n3558), .Y(n2881) );
  OAI21X1 U2617 ( .A(n5733), .B(n5780), .C(n4061), .Y(n2882) );
  OAI21X1 U2619 ( .A(n5732), .B(n5781), .C(n4147), .Y(n2883) );
  OAI21X1 U2621 ( .A(n5731), .B(n5780), .C(n4237), .Y(n2884) );
  OAI21X1 U2623 ( .A(n5749), .B(n5781), .C(n3320), .Y(n2885) );
  OAI21X1 U2625 ( .A(n5750), .B(n5780), .C(n3635), .Y(n2886) );
  OAI21X1 U2627 ( .A(n5751), .B(n5780), .C(n3718), .Y(n2887) );
  OAI21X1 U2629 ( .A(n5752), .B(n5781), .C(n3801), .Y(n2888) );
  OAI21X1 U2631 ( .A(n5753), .B(n5780), .C(n3885), .Y(n2889) );
  OAI21X1 U2633 ( .A(n5754), .B(n5780), .C(n3969), .Y(n2890) );
  OAI21X1 U2635 ( .A(n5755), .B(n5781), .C(n3399), .Y(n2891) );
  OAI21X1 U2637 ( .A(n5756), .B(n5781), .C(n3478), .Y(n2892) );
  OAI21X1 U2639 ( .A(n5757), .B(n5780), .C(n3557), .Y(n2893) );
  OAI21X1 U2641 ( .A(n5758), .B(n5781), .C(n4060), .Y(n2894) );
  OAI21X1 U2643 ( .A(n5759), .B(n5780), .C(n4146), .Y(n2895) );
  OAI21X1 U2645 ( .A(n5760), .B(n5780), .C(n3717), .Y(n2896) );
  OAI21X1 U2647 ( .A(n5761), .B(n5781), .C(n3800), .Y(n2897) );
  OAI21X1 U2649 ( .A(n5762), .B(n5781), .C(n3884), .Y(n2898) );
  OAI21X1 U2651 ( .A(n5763), .B(n5781), .C(n3556), .Y(n2899) );
  OAI21X1 U2653 ( .A(n5764), .B(n5780), .C(n3020), .Y(n2900) );
  OAI21X1 U2655 ( .A(n5765), .B(n5781), .C(n3095), .Y(n2901) );
  OAI21X1 U2657 ( .A(n5766), .B(n5781), .C(n3170), .Y(n2902) );
  OAI21X1 U2659 ( .A(n5767), .B(n5781), .C(n3247), .Y(n2903) );
  OAI21X1 U2661 ( .A(n5768), .B(n5780), .C(n120), .Y(n2904) );
  OAI21X1 U2663 ( .A(n5769), .B(n5781), .C(n3398), .Y(n2905) );
  OAI21X1 U2665 ( .A(n5770), .B(n5780), .C(n3019), .Y(n2906) );
  OAI21X1 U2667 ( .A(n5771), .B(n5781), .C(n3094), .Y(n2907) );
  OAI21X1 U2669 ( .A(n5772), .B(n5780), .C(n3477), .Y(n2908) );
  OAI21X1 U2671 ( .A(n5748), .B(n5781), .C(n3246), .Y(n2909) );
  OAI21X1 U2673 ( .A(n5747), .B(n5780), .C(n119), .Y(n2910) );
  NOR3X1 U2676 ( .A(n5898), .B(wr_ptr[1]), .C(n5900), .Y(n442) );
  OAI21X1 U2677 ( .A(n5746), .B(n5778), .C(n3883), .Y(n2911) );
  OAI21X1 U2679 ( .A(n5745), .B(n5778), .C(n3799), .Y(n2912) );
  OAI21X1 U2681 ( .A(n5744), .B(n5778), .C(n3716), .Y(n2913) );
  OAI21X1 U2683 ( .A(n5743), .B(n5779), .C(n3634), .Y(n2914) );
  OAI21X1 U2685 ( .A(n5742), .B(n5778), .C(n4236), .Y(n2915) );
  OAI21X1 U2687 ( .A(n5741), .B(n5779), .C(n4145), .Y(n2916) );
  OAI21X1 U2689 ( .A(n5740), .B(n5779), .C(n4059), .Y(n2917) );
  OAI21X1 U2691 ( .A(n5739), .B(n5779), .C(n3968), .Y(n2918) );
  OAI21X1 U2693 ( .A(n5738), .B(n5778), .C(n3882), .Y(n2919) );
  OAI21X1 U2695 ( .A(n5737), .B(n5778), .C(n3245), .Y(n2920) );
  OAI21X1 U2697 ( .A(n5736), .B(n5779), .C(n3169), .Y(n2921) );
  OAI21X1 U2699 ( .A(n5735), .B(n5778), .C(n3093), .Y(n2922) );
  OAI21X1 U2701 ( .A(n5734), .B(n5779), .C(n3018), .Y(n2923) );
  OAI21X1 U2703 ( .A(n5733), .B(n5778), .C(n3798), .Y(n2924) );
  OAI21X1 U2705 ( .A(n5732), .B(n5779), .C(n3715), .Y(n2925) );
  OAI21X1 U2707 ( .A(n5731), .B(n5778), .C(n3633), .Y(n2926) );
  OAI21X1 U2709 ( .A(n5749), .B(n5779), .C(n3244), .Y(n2927) );
  OAI21X1 U2711 ( .A(n5750), .B(n5778), .C(n4235), .Y(n2928) );
  OAI21X1 U2713 ( .A(n5751), .B(n5778), .C(n4144), .Y(n2929) );
  OAI21X1 U2715 ( .A(n5752), .B(n5779), .C(n4058), .Y(n2930) );
  OAI21X1 U2717 ( .A(n5753), .B(n5778), .C(n3967), .Y(n2931) );
  OAI21X1 U2719 ( .A(n5754), .B(n5778), .C(n3881), .Y(n2932) );
  OAI21X1 U2721 ( .A(n5755), .B(n5779), .C(n3168), .Y(n2933) );
  OAI21X1 U2723 ( .A(n5756), .B(n5779), .C(n3092), .Y(n2934) );
  OAI21X1 U2725 ( .A(n5757), .B(n5778), .C(n3017), .Y(n2935) );
  OAI21X1 U2727 ( .A(n5758), .B(n5779), .C(n3797), .Y(n2936) );
  OAI21X1 U2729 ( .A(n5759), .B(n5778), .C(n3714), .Y(n2937) );
  OAI21X1 U2731 ( .A(n5760), .B(n5778), .C(n4143), .Y(n2938) );
  OAI21X1 U2733 ( .A(n5761), .B(n5779), .C(n4057), .Y(n2939) );
  OAI21X1 U2735 ( .A(n5762), .B(n5779), .C(n3966), .Y(n2940) );
  OAI21X1 U2737 ( .A(n5763), .B(n5779), .C(n3016), .Y(n2941) );
  OAI21X1 U2739 ( .A(n5764), .B(n5778), .C(n3555), .Y(n2942) );
  OAI21X1 U2741 ( .A(n5765), .B(n5779), .C(n3476), .Y(n2943) );
  OAI21X1 U2743 ( .A(n5766), .B(n5779), .C(n3397), .Y(n2944) );
  OAI21X1 U2745 ( .A(n5767), .B(n5779), .C(n3319), .Y(n2945) );
  OAI21X1 U2747 ( .A(n5768), .B(n5778), .C(n118), .Y(n2946) );
  OAI21X1 U2749 ( .A(n5769), .B(n5779), .C(n3167), .Y(n2947) );
  OAI21X1 U2751 ( .A(n5770), .B(n5778), .C(n3554), .Y(n2948) );
  OAI21X1 U2753 ( .A(n5771), .B(n5779), .C(n3475), .Y(n2949) );
  OAI21X1 U2755 ( .A(n5772), .B(n5778), .C(n3091), .Y(n2950) );
  OAI21X1 U2757 ( .A(n5748), .B(n5779), .C(n3318), .Y(n2951) );
  OAI21X1 U2759 ( .A(n5747), .B(n5778), .C(n117), .Y(n2952) );
  NOR3X1 U2762 ( .A(n5899), .B(wr_ptr[0]), .C(n5900), .Y(n486) );
  OAI21X1 U2763 ( .A(n5746), .B(n5776), .C(n3796), .Y(n2953) );
  OAI21X1 U2765 ( .A(n5745), .B(n5776), .C(n3880), .Y(n2954) );
  OAI21X1 U2767 ( .A(n5744), .B(n5776), .C(n3632), .Y(n2955) );
  OAI21X1 U2769 ( .A(n5743), .B(n5777), .C(n3713), .Y(n2956) );
  OAI21X1 U2771 ( .A(n5742), .B(n5776), .C(n4142), .Y(n2957) );
  OAI21X1 U2773 ( .A(n5741), .B(n5777), .C(n4234), .Y(n2958) );
  OAI21X1 U2775 ( .A(n5740), .B(n5777), .C(n3965), .Y(n2959) );
  OAI21X1 U2777 ( .A(n5739), .B(n5777), .C(n4056), .Y(n2960) );
  OAI21X1 U2779 ( .A(n5738), .B(n5776), .C(n3795), .Y(n2961) );
  OAI21X1 U2781 ( .A(n5737), .B(n5776), .C(n3166), .Y(n2962) );
  OAI21X1 U2783 ( .A(n5736), .B(n5777), .C(n3243), .Y(n2963) );
  OAI21X1 U2785 ( .A(n5735), .B(n5776), .C(n3015), .Y(n2964) );
  OAI21X1 U2787 ( .A(n5734), .B(n5777), .C(n3090), .Y(n2965) );
  OAI21X1 U2789 ( .A(n5733), .B(n5776), .C(n3879), .Y(n2966) );
  OAI21X1 U2791 ( .A(n5732), .B(n5777), .C(n3631), .Y(n2967) );
  OAI21X1 U2793 ( .A(n5731), .B(n5776), .C(n3712), .Y(n2968) );
  OAI21X1 U2795 ( .A(n5749), .B(n5777), .C(n3165), .Y(n2969) );
  OAI21X1 U2797 ( .A(n5750), .B(n5776), .C(n4141), .Y(n2970) );
  OAI21X1 U2799 ( .A(n5751), .B(n5776), .C(n4233), .Y(n2971) );
  OAI21X1 U2801 ( .A(n5752), .B(n5777), .C(n3964), .Y(n2972) );
  OAI21X1 U2803 ( .A(n5753), .B(n5776), .C(n4055), .Y(n2973) );
  OAI21X1 U2805 ( .A(n5754), .B(n5776), .C(n3794), .Y(n2974) );
  OAI21X1 U2807 ( .A(n5755), .B(n5777), .C(n3242), .Y(n2975) );
  OAI21X1 U2809 ( .A(n5756), .B(n5777), .C(n3014), .Y(n2976) );
  OAI21X1 U2811 ( .A(n5757), .B(n5776), .C(n3089), .Y(n2977) );
  OAI21X1 U2813 ( .A(n5758), .B(n5777), .C(n3878), .Y(n2978) );
  OAI21X1 U2815 ( .A(n5759), .B(n5776), .C(n3630), .Y(n2979) );
  OAI21X1 U2817 ( .A(n5760), .B(n5776), .C(n4232), .Y(n2980) );
  OAI21X1 U2819 ( .A(n5761), .B(n5777), .C(n3963), .Y(n2981) );
  OAI21X1 U2821 ( .A(n5762), .B(n5777), .C(n4054), .Y(n2982) );
  OAI21X1 U2823 ( .A(n5763), .B(n5777), .C(n3088), .Y(n2983) );
  OAI21X1 U2825 ( .A(n5764), .B(n5776), .C(n3474), .Y(n2984) );
  OAI21X1 U2827 ( .A(n5765), .B(n5777), .C(n3553), .Y(n2985) );
  OAI21X1 U2829 ( .A(n5766), .B(n5777), .C(n3317), .Y(n2986) );
  OAI21X1 U2831 ( .A(n5767), .B(n5777), .C(n3396), .Y(n2987) );
  OAI21X1 U2833 ( .A(n5768), .B(n5776), .C(n116), .Y(n2988) );
  OAI21X1 U2835 ( .A(n5769), .B(n5777), .C(n3241), .Y(n2989) );
  OAI21X1 U2837 ( .A(n5770), .B(n5776), .C(n3473), .Y(n2990) );
  OAI21X1 U2839 ( .A(n5771), .B(n5777), .C(n3552), .Y(n2991) );
  OAI21X1 U2841 ( .A(n5772), .B(n5776), .C(n3013), .Y(n2992) );
  OAI21X1 U2843 ( .A(n5748), .B(n5777), .C(n3395), .Y(n2993) );
  OAI21X1 U2845 ( .A(n5747), .B(n5776), .C(n115), .Y(n2994) );
  NOR3X1 U2848 ( .A(n5899), .B(n5898), .C(n5900), .Y(n530) );
  NOR3X1 U2849 ( .A(n5901), .B(n1568), .C(n5902), .Y(n1264) );
  OAI21X1 U2850 ( .A(n5902), .B(n4322), .C(n3961), .Y(n2995) );
  OAI21X1 U2852 ( .A(n5901), .B(n4322), .C(n3876), .Y(n2996) );
  OAI21X1 U2854 ( .A(n5900), .B(n4322), .C(n3792), .Y(n2997) );
  OAI21X1 U2856 ( .A(n5899), .B(n4322), .C(n3710), .Y(n2998) );
  OAI21X1 U2858 ( .A(n5898), .B(n4322), .C(n3629), .Y(n2999) );
  OAI21X1 U2862 ( .A(n1575), .B(n5903), .C(n114), .Y(n3000) );
  AOI22X1 U2863 ( .A(n107), .B(n1577), .C(n95), .D(n1578), .Y(n1576) );
  OAI21X1 U2864 ( .A(n1575), .B(n5850), .C(n113), .Y(n3001) );
  AOI22X1 U2865 ( .A(n106), .B(n1577), .C(n94), .D(n1578), .Y(n1579) );
  OAI21X1 U2866 ( .A(n1575), .B(n5851), .C(n112), .Y(n3002) );
  AOI22X1 U2867 ( .A(n105), .B(n1577), .C(n93), .D(n1578), .Y(n1580) );
  OAI21X1 U2868 ( .A(n1575), .B(n5904), .C(n111), .Y(n3003) );
  AOI22X1 U2869 ( .A(n104), .B(n1577), .C(n92), .D(n1578), .Y(n1581) );
  OAI21X1 U2870 ( .A(n1575), .B(n103), .C(n110), .Y(n3004) );
  AOI22X1 U2871 ( .A(n103), .B(n1577), .C(n103), .D(n1578), .Y(n1582) );
  OAI21X1 U2872 ( .A(n4230), .B(n5840), .C(n4053), .Y(n3005) );
  OAI21X1 U2874 ( .A(n4230), .B(n5841), .C(n3962), .Y(n3006) );
  OAI21X1 U2876 ( .A(n4230), .B(n5842), .C(n3877), .Y(n3007) );
  OAI21X1 U2878 ( .A(n4230), .B(n5843), .C(n3793), .Y(n3008) );
  OAI21X1 U2880 ( .A(n4230), .B(n5844), .C(n3711), .Y(n3009) );
  AOI22X1 U2883 ( .A(data_out[41]), .B(n4323), .C(n24), .D(n5775), .Y(n1590)
         );
  AOI22X1 U2884 ( .A(data_out[40]), .B(n4323), .C(n25), .D(n5773), .Y(n1591)
         );
  AOI22X1 U2885 ( .A(data_out[39]), .B(n4323), .C(n26), .D(n5773), .Y(n1592)
         );
  AOI22X1 U2886 ( .A(data_out[38]), .B(n4323), .C(n27), .D(n5773), .Y(n1593)
         );
  AOI22X1 U2887 ( .A(data_out[37]), .B(n4323), .C(n28), .D(n5773), .Y(n1594)
         );
  AOI22X1 U2888 ( .A(data_out[36]), .B(n4323), .C(n29), .D(n5773), .Y(n1595)
         );
  AOI22X1 U2889 ( .A(data_out[35]), .B(n4323), .C(n30), .D(n5775), .Y(n1596)
         );
  AOI22X1 U2890 ( .A(data_out[34]), .B(n4323), .C(n31), .D(n5773), .Y(n1597)
         );
  AOI22X1 U2891 ( .A(data_out[33]), .B(n4323), .C(n32), .D(n5773), .Y(n1598)
         );
  AOI22X1 U2892 ( .A(data_out[32]), .B(n4323), .C(n33), .D(n5775), .Y(n1599)
         );
  AOI22X1 U2893 ( .A(data_out[31]), .B(n4323), .C(n34), .D(n5773), .Y(n1600)
         );
  AOI22X1 U2894 ( .A(data_out[30]), .B(n5774), .C(n35), .D(n5775), .Y(n1601)
         );
  AOI22X1 U2895 ( .A(data_out[29]), .B(n5774), .C(n36), .D(n5773), .Y(n1602)
         );
  AOI22X1 U2896 ( .A(data_out[28]), .B(n5774), .C(n37), .D(n5773), .Y(n1603)
         );
  AOI22X1 U2897 ( .A(data_out[27]), .B(n5774), .C(n38), .D(n5775), .Y(n1604)
         );
  AOI22X1 U2898 ( .A(data_out[26]), .B(n5774), .C(n39), .D(n5773), .Y(n1605)
         );
  AOI22X1 U2899 ( .A(data_out[25]), .B(n5774), .C(n40), .D(n5775), .Y(n1606)
         );
  AOI22X1 U2900 ( .A(data_out[24]), .B(n5774), .C(n41), .D(n5773), .Y(n1607)
         );
  AOI22X1 U2901 ( .A(data_out[23]), .B(n5774), .C(n42), .D(n5773), .Y(n1608)
         );
  AOI22X1 U2902 ( .A(data_out[22]), .B(n5774), .C(n43), .D(n5773), .Y(n1609)
         );
  AOI22X1 U2903 ( .A(data_out[21]), .B(n5774), .C(n44), .D(n5773), .Y(n1610)
         );
  AOI22X1 U2904 ( .A(data_out[20]), .B(n5774), .C(n45), .D(n5773), .Y(n1611)
         );
  AOI22X1 U2905 ( .A(data_out[19]), .B(n5774), .C(n46), .D(n5773), .Y(n1612)
         );
  AOI22X1 U2906 ( .A(data_out[18]), .B(n5774), .C(n47), .D(n5773), .Y(n1613)
         );
  AOI22X1 U2907 ( .A(data_out[17]), .B(n5774), .C(n48), .D(n5773), .Y(n1614)
         );
  AOI22X1 U2908 ( .A(data_out[16]), .B(n5774), .C(n49), .D(n5773), .Y(n1615)
         );
  AOI22X1 U2909 ( .A(data_out[15]), .B(n5774), .C(n50), .D(n5773), .Y(n1616)
         );
  AOI22X1 U2910 ( .A(data_out[14]), .B(n5774), .C(n51), .D(n5773), .Y(n1617)
         );
  AOI22X1 U2911 ( .A(data_out[13]), .B(n5774), .C(n52), .D(n5773), .Y(n1618)
         );
  AOI22X1 U2912 ( .A(data_out[12]), .B(n5774), .C(n53), .D(n5773), .Y(n1619)
         );
  AOI22X1 U2913 ( .A(data_out[11]), .B(n5774), .C(n54), .D(n5773), .Y(n1620)
         );
  AOI22X1 U2914 ( .A(data_out[10]), .B(n5774), .C(n55), .D(n5773), .Y(n1621)
         );
  AOI22X1 U2915 ( .A(data_out[9]), .B(n5774), .C(n56), .D(n5775), .Y(n1622) );
  AOI22X1 U2916 ( .A(data_out[8]), .B(n5774), .C(n57), .D(n5773), .Y(n1623) );
  AOI22X1 U2917 ( .A(data_out[7]), .B(n5774), .C(n58), .D(n5773), .Y(n1624) );
  AOI22X1 U2918 ( .A(data_out[6]), .B(n5774), .C(n59), .D(n5773), .Y(n1625) );
  AOI22X1 U2919 ( .A(data_out[5]), .B(n5774), .C(n60), .D(n5773), .Y(n1626) );
  AOI22X1 U2920 ( .A(data_out[4]), .B(n5774), .C(n61), .D(n5773), .Y(n1627) );
  AOI22X1 U2921 ( .A(data_out[3]), .B(n5774), .C(n62), .D(n5775), .Y(n1628) );
  AOI22X1 U2922 ( .A(data_out[2]), .B(n5774), .C(n63), .D(n5773), .Y(n1629) );
  AOI22X1 U2923 ( .A(data_out[1]), .B(n5774), .C(n64), .D(n5773), .Y(n1630) );
  AOI22X1 U2924 ( .A(data_out[0]), .B(n5774), .C(n65), .D(n5773), .Y(n1631) );
  OAI21X1 U2926 ( .A(n4051), .B(n5897), .C(n4050), .Y(n3010) );
  NAND3X1 U2928 ( .A(n4052), .B(n5845), .C(n4140), .Y(n1634) );
  NAND3X1 U2929 ( .A(n1638), .B(n5894), .C(n1639), .Y(n1637) );
  NOR3X1 U2930 ( .A(n4318), .B(fillcount[3]), .C(fillcount[2]), .Y(n1639) );
  OAI21X1 U2932 ( .A(n1575), .B(n5896), .C(n109), .Y(n3011) );
  AOI22X1 U2933 ( .A(n108), .B(n1577), .C(n96), .D(n1578), .Y(n1641) );
  OAI21X1 U2935 ( .A(n3959), .B(n5895), .C(n3958), .Y(n3012) );
  NAND3X1 U2937 ( .A(n3960), .B(n5845), .C(n4321), .Y(n1644) );
  NAND3X1 U2938 ( .A(get), .B(n5897), .C(n1643), .Y(n1632) );
  NAND3X1 U2939 ( .A(n4139), .B(n1573), .C(n1649), .Y(n1646) );
  NOR3X1 U2940 ( .A(n4227), .B(fillcount[5]), .C(n5903), .Y(n1649) );
  NAND3X1 U2943 ( .A(n1647), .B(n5897), .C(get), .Y(n1633) );
  HAX1 add_45_U1_1_1 ( .A(fillcount[1]), .B(fillcount[0]), .YC(add_45_carry[2]), .YS(n92) );
  HAX1 add_45_U1_1_2 ( .A(fillcount[2]), .B(add_45_carry[2]), .YC(
        add_45_carry[3]), .YS(n93) );
  HAX1 add_45_U1_1_3 ( .A(fillcount[3]), .B(add_45_carry[3]), .YC(
        add_45_carry[4]), .YS(n94) );
  HAX1 add_45_U1_1_4 ( .A(fillcount[4]), .B(add_45_carry[4]), .YC(
        add_45_carry[5]), .YS(n95) );
  HAX1 r308_U1_1_1 ( .A(n5706), .B(n5646), .YC(r308_carry[2]), .YS(n81) );
  HAX1 r308_U1_1_2 ( .A(n5730), .B(r308_carry[2]), .YC(r308_carry[3]), .YS(n82) );
  HAX1 r308_U1_1_3 ( .A(n22), .B(r308_carry[3]), .YC(r308_carry[4]), .YS(n83)
         );
  HAX1 r307_U1_1_1 ( .A(wr_ptr[1]), .B(wr_ptr[0]), .YC(r307_carry[2]), .YS(n76) );
  HAX1 r307_U1_1_2 ( .A(wr_ptr[2]), .B(r307_carry[2]), .YC(r307_carry[3]), 
        .YS(n77) );
  HAX1 r307_U1_1_3 ( .A(wr_ptr[3]), .B(r307_carry[3]), .YC(r307_carry[4]), 
        .YS(n78) );
  OR2X1 U3 ( .A(n3957), .B(reset), .Y(n1574) );
  OR2X1 U4 ( .A(n3875), .B(n1573), .Y(n1575) );
  OR2X1 U5 ( .A(n4320), .B(fillcount[4]), .Y(n5849) );
  AND2X1 U6 ( .A(n4051), .B(n3875), .Y(n1635) );
  AND2X1 U7 ( .A(n1573), .B(n3959), .Y(n1645) );
  AND2X1 U8 ( .A(n1574), .B(n4321), .Y(n4323) );
  AND2X1 U9 ( .A(n4140), .B(n1574), .Y(n1568) );
  AND2X1 U10 ( .A(n1642), .B(n3957), .Y(n1573) );
  BUFX2 U11 ( .A(n1631), .Y(n1) );
  BUFX2 U12 ( .A(n1630), .Y(n2) );
  BUFX2 U13 ( .A(n1629), .Y(n3) );
  BUFX2 U14 ( .A(n1628), .Y(n4) );
  BUFX2 U15 ( .A(n1627), .Y(n5) );
  BUFX2 U16 ( .A(n1626), .Y(n6) );
  BUFX2 U17 ( .A(n1625), .Y(n7) );
  BUFX2 U18 ( .A(n1624), .Y(n8) );
  BUFX2 U19 ( .A(n1623), .Y(n9) );
  BUFX2 U20 ( .A(n1622), .Y(n10) );
  BUFX2 U21 ( .A(n1621), .Y(n11) );
  BUFX2 U22 ( .A(n1620), .Y(n12) );
  BUFX2 U23 ( .A(n1619), .Y(n13) );
  BUFX2 U24 ( .A(n1618), .Y(n14) );
  BUFX2 U25 ( .A(n1617), .Y(n15) );
  BUFX2 U26 ( .A(n1616), .Y(n16) );
  BUFX2 U27 ( .A(n1615), .Y(n17) );
  BUFX2 U28 ( .A(n1614), .Y(n18) );
  BUFX2 U29 ( .A(n1613), .Y(n66) );
  BUFX2 U30 ( .A(n1612), .Y(n67) );
  BUFX2 U31 ( .A(n1611), .Y(n68) );
  BUFX2 U32 ( .A(n1610), .Y(n69) );
  BUFX2 U33 ( .A(n1609), .Y(n70) );
  BUFX2 U34 ( .A(n1608), .Y(n71) );
  BUFX2 U35 ( .A(n1607), .Y(n72) );
  BUFX2 U36 ( .A(n1606), .Y(n73) );
  BUFX2 U37 ( .A(n1605), .Y(n74) );
  BUFX2 U38 ( .A(n1604), .Y(n75) );
  BUFX2 U39 ( .A(n1603), .Y(n80) );
  BUFX2 U40 ( .A(n1602), .Y(n85) );
  BUFX2 U41 ( .A(n1601), .Y(n86) );
  BUFX2 U42 ( .A(n1600), .Y(n87) );
  BUFX2 U43 ( .A(n1599), .Y(n88) );
  BUFX2 U44 ( .A(n1598), .Y(n89) );
  BUFX2 U45 ( .A(n1597), .Y(n90) );
  BUFX2 U46 ( .A(n1596), .Y(n91) );
  BUFX2 U47 ( .A(n1595), .Y(n97) );
  BUFX2 U48 ( .A(n1594), .Y(n98) );
  BUFX2 U49 ( .A(n1593), .Y(n99) );
  BUFX2 U50 ( .A(n1592), .Y(n100) );
  BUFX2 U51 ( .A(n1591), .Y(n101) );
  BUFX2 U52 ( .A(n1590), .Y(n102) );
  AND2X1 U53 ( .A(n1264), .B(n530), .Y(n1523) );
  AND2X1 U54 ( .A(n1264), .B(n486), .Y(n1480) );
  AND2X1 U55 ( .A(n1264), .B(n442), .Y(n1437) );
  AND2X1 U56 ( .A(n1264), .B(n398), .Y(n1394) );
  AND2X1 U57 ( .A(n1264), .B(n354), .Y(n1351) );
  AND2X1 U58 ( .A(n1264), .B(n310), .Y(n1308) );
  AND2X1 U59 ( .A(n1264), .B(n266), .Y(n1265) );
  AND2X1 U60 ( .A(n1264), .B(n221), .Y(n1221) );
  AND2X1 U61 ( .A(n919), .B(n530), .Y(n1178) );
  AND2X1 U62 ( .A(n919), .B(n486), .Y(n1135) );
  AND2X1 U63 ( .A(n919), .B(n442), .Y(n1092) );
  AND2X1 U64 ( .A(n919), .B(n398), .Y(n1049) );
  AND2X1 U65 ( .A(n919), .B(n354), .Y(n1006) );
  AND2X1 U66 ( .A(n919), .B(n310), .Y(n963) );
  AND2X1 U67 ( .A(n919), .B(n266), .Y(n920) );
  AND2X1 U68 ( .A(n919), .B(n221), .Y(n876) );
  AND2X1 U69 ( .A(n574), .B(n530), .Y(n833) );
  AND2X1 U70 ( .A(n574), .B(n486), .Y(n790) );
  AND2X1 U71 ( .A(n574), .B(n442), .Y(n747) );
  AND2X1 U72 ( .A(n574), .B(n398), .Y(n704) );
  AND2X1 U73 ( .A(n574), .B(n354), .Y(n661) );
  AND2X1 U74 ( .A(n574), .B(n310), .Y(n618) );
  AND2X1 U75 ( .A(n574), .B(n266), .Y(n575) );
  AND2X1 U76 ( .A(n574), .B(n221), .Y(n531) );
  AND2X1 U77 ( .A(n530), .B(n222), .Y(n487) );
  AND2X1 U78 ( .A(n486), .B(n222), .Y(n443) );
  AND2X1 U79 ( .A(n442), .B(n222), .Y(n399) );
  AND2X1 U80 ( .A(n398), .B(n222), .Y(n355) );
  AND2X1 U81 ( .A(n354), .B(n222), .Y(n311) );
  AND2X1 U82 ( .A(n310), .B(n222), .Y(n267) );
  AND2X1 U83 ( .A(n266), .B(n222), .Y(n223) );
  AND2X1 U84 ( .A(n221), .B(n222), .Y(n178) );
  BUFX2 U85 ( .A(n1641), .Y(n109) );
  BUFX2 U86 ( .A(n1582), .Y(n110) );
  BUFX2 U87 ( .A(n1581), .Y(n111) );
  BUFX2 U88 ( .A(n1580), .Y(n112) );
  BUFX2 U89 ( .A(n1579), .Y(n113) );
  BUFX2 U90 ( .A(n1576), .Y(n114) );
  AND2X1 U91 ( .A(fifo_array[1343]), .B(n5777), .Y(n1565) );
  INVX1 U92 ( .A(n1565), .Y(n115) );
  AND2X1 U93 ( .A(fifo_array[1337]), .B(n5776), .Y(n1559) );
  INVX1 U94 ( .A(n1559), .Y(n116) );
  AND2X1 U95 ( .A(fifo_array[1301]), .B(n5779), .Y(n1522) );
  INVX1 U96 ( .A(n1522), .Y(n117) );
  AND2X1 U97 ( .A(fifo_array[1295]), .B(n5778), .Y(n1516) );
  INVX1 U98 ( .A(n1516), .Y(n118) );
  AND2X1 U99 ( .A(fifo_array[1259]), .B(n5781), .Y(n1479) );
  INVX1 U100 ( .A(n1479), .Y(n119) );
  AND2X1 U101 ( .A(fifo_array[1253]), .B(n5780), .Y(n1473) );
  INVX1 U102 ( .A(n1473), .Y(n120) );
  AND2X1 U103 ( .A(fifo_array[1217]), .B(n5783), .Y(n1436) );
  INVX1 U104 ( .A(n1436), .Y(n121) );
  AND2X1 U105 ( .A(fifo_array[1211]), .B(n5782), .Y(n1430) );
  INVX1 U106 ( .A(n1430), .Y(n122) );
  AND2X1 U107 ( .A(fifo_array[1175]), .B(n5785), .Y(n1393) );
  INVX1 U108 ( .A(n1393), .Y(n123) );
  AND2X1 U109 ( .A(fifo_array[1169]), .B(n5784), .Y(n1387) );
  INVX1 U110 ( .A(n1387), .Y(n124) );
  AND2X1 U111 ( .A(fifo_array[1133]), .B(n5787), .Y(n1350) );
  INVX1 U112 ( .A(n1350), .Y(n125) );
  AND2X1 U113 ( .A(fifo_array[1127]), .B(n5786), .Y(n1344) );
  INVX1 U114 ( .A(n1344), .Y(n126) );
  AND2X1 U115 ( .A(fifo_array[1091]), .B(n5789), .Y(n1307) );
  INVX1 U116 ( .A(n1307), .Y(n127) );
  AND2X1 U117 ( .A(fifo_array[1085]), .B(n5789), .Y(n1301) );
  INVX1 U119 ( .A(n1301), .Y(n128) );
  AND2X1 U121 ( .A(fifo_array[1049]), .B(n5791), .Y(n1263) );
  INVX1 U123 ( .A(n1263), .Y(n129) );
  AND2X1 U125 ( .A(fifo_array[1043]), .B(n5791), .Y(n1257) );
  INVX1 U127 ( .A(n1257), .Y(n130) );
  AND2X1 U129 ( .A(fifo_array[1007]), .B(n5792), .Y(n1220) );
  INVX1 U131 ( .A(n1220), .Y(n131) );
  AND2X1 U133 ( .A(fifo_array[1001]), .B(n5793), .Y(n1214) );
  INVX1 U135 ( .A(n1214), .Y(n132) );
  AND2X1 U137 ( .A(fifo_array[965]), .B(n5794), .Y(n1177) );
  INVX1 U139 ( .A(n1177), .Y(n133) );
  AND2X1 U141 ( .A(fifo_array[959]), .B(n5795), .Y(n1171) );
  INVX1 U143 ( .A(n1171), .Y(n134) );
  AND2X1 U145 ( .A(fifo_array[923]), .B(n5796), .Y(n1134) );
  INVX1 U147 ( .A(n1134), .Y(n135) );
  AND2X1 U149 ( .A(fifo_array[917]), .B(n5797), .Y(n1128) );
  INVX1 U151 ( .A(n1128), .Y(n136) );
  AND2X1 U153 ( .A(fifo_array[881]), .B(n5798), .Y(n1091) );
  INVX1 U155 ( .A(n1091), .Y(n137) );
  AND2X1 U157 ( .A(fifo_array[875]), .B(n5799), .Y(n1085) );
  INVX1 U159 ( .A(n1085), .Y(n138) );
  AND2X1 U161 ( .A(fifo_array[839]), .B(n5800), .Y(n1048) );
  INVX1 U163 ( .A(n1048), .Y(n139) );
  AND2X1 U165 ( .A(fifo_array[833]), .B(n5801), .Y(n1042) );
  INVX1 U167 ( .A(n1042), .Y(n140) );
  AND2X1 U169 ( .A(fifo_array[797]), .B(n5802), .Y(n1005) );
  INVX1 U171 ( .A(n1005), .Y(n141) );
  AND2X1 U173 ( .A(fifo_array[791]), .B(n5803), .Y(n999) );
  INVX1 U175 ( .A(n999), .Y(n142) );
  AND2X1 U177 ( .A(fifo_array[755]), .B(n5804), .Y(n962) );
  INVX1 U179 ( .A(n962), .Y(n143) );
  AND2X1 U181 ( .A(fifo_array[749]), .B(n5805), .Y(n956) );
  INVX1 U183 ( .A(n956), .Y(n144) );
  AND2X1 U185 ( .A(fifo_array[713]), .B(n5806), .Y(n918) );
  INVX1 U187 ( .A(n918), .Y(n145) );
  AND2X1 U189 ( .A(fifo_array[707]), .B(n5807), .Y(n912) );
  INVX1 U191 ( .A(n912), .Y(n146) );
  AND2X1 U193 ( .A(fifo_array[671]), .B(n5808), .Y(n875) );
  INVX1 U195 ( .A(n875), .Y(n147) );
  AND2X1 U197 ( .A(fifo_array[665]), .B(n5809), .Y(n869) );
  INVX1 U199 ( .A(n869), .Y(n148) );
  AND2X1 U201 ( .A(fifo_array[629]), .B(n5810), .Y(n832) );
  INVX1 U202 ( .A(n832), .Y(n149) );
  AND2X1 U204 ( .A(fifo_array[623]), .B(n5811), .Y(n826) );
  INVX1 U206 ( .A(n826), .Y(n150) );
  AND2X1 U208 ( .A(fifo_array[587]), .B(n5812), .Y(n789) );
  INVX1 U210 ( .A(n789), .Y(n151) );
  AND2X1 U212 ( .A(fifo_array[581]), .B(n5813), .Y(n783) );
  INVX1 U214 ( .A(n783), .Y(n152) );
  AND2X1 U216 ( .A(fifo_array[545]), .B(n5814), .Y(n746) );
  INVX1 U218 ( .A(n746), .Y(n153) );
  AND2X1 U220 ( .A(fifo_array[539]), .B(n5815), .Y(n740) );
  INVX1 U222 ( .A(n740), .Y(n154) );
  AND2X1 U224 ( .A(fifo_array[503]), .B(n5816), .Y(n703) );
  INVX1 U226 ( .A(n703), .Y(n155) );
  AND2X1 U228 ( .A(fifo_array[497]), .B(n5817), .Y(n697) );
  INVX1 U230 ( .A(n697), .Y(n156) );
  AND2X1 U232 ( .A(fifo_array[461]), .B(n5818), .Y(n660) );
  INVX1 U234 ( .A(n660), .Y(n157) );
  AND2X1 U236 ( .A(fifo_array[455]), .B(n5819), .Y(n654) );
  INVX1 U238 ( .A(n654), .Y(n158) );
  AND2X1 U240 ( .A(fifo_array[419]), .B(n5820), .Y(n617) );
  INVX1 U242 ( .A(n617), .Y(n159) );
  AND2X1 U244 ( .A(fifo_array[413]), .B(n5821), .Y(n611) );
  INVX1 U246 ( .A(n611), .Y(n160) );
  AND2X1 U248 ( .A(fifo_array[377]), .B(n5822), .Y(n573) );
  INVX1 U250 ( .A(n573), .Y(n161) );
  AND2X1 U252 ( .A(fifo_array[371]), .B(n5823), .Y(n567) );
  INVX1 U254 ( .A(n567), .Y(n162) );
  AND2X1 U256 ( .A(fifo_array[335]), .B(n5824), .Y(n529) );
  INVX1 U258 ( .A(n529), .Y(n163) );
  AND2X1 U260 ( .A(fifo_array[329]), .B(n5825), .Y(n523) );
  INVX1 U262 ( .A(n523), .Y(n164) );
  AND2X1 U264 ( .A(fifo_array[293]), .B(n5826), .Y(n485) );
  INVX1 U266 ( .A(n485), .Y(n165) );
  AND2X1 U268 ( .A(fifo_array[287]), .B(n5827), .Y(n479) );
  INVX1 U270 ( .A(n479), .Y(n166) );
  AND2X1 U272 ( .A(fifo_array[251]), .B(n5828), .Y(n441) );
  INVX1 U274 ( .A(n441), .Y(n167) );
  AND2X1 U276 ( .A(fifo_array[245]), .B(n5829), .Y(n435) );
  INVX1 U278 ( .A(n435), .Y(n168) );
  AND2X1 U280 ( .A(fifo_array[209]), .B(n5830), .Y(n397) );
  INVX1 U282 ( .A(n397), .Y(n169) );
  AND2X1 U284 ( .A(fifo_array[203]), .B(n5831), .Y(n391) );
  INVX1 U286 ( .A(n391), .Y(n170) );
  AND2X1 U287 ( .A(fifo_array[167]), .B(n5832), .Y(n353) );
  INVX1 U289 ( .A(n353), .Y(n171) );
  AND2X1 U291 ( .A(fifo_array[161]), .B(n5833), .Y(n347) );
  INVX1 U293 ( .A(n347), .Y(n172) );
  AND2X1 U295 ( .A(fifo_array[125]), .B(n5834), .Y(n309) );
  INVX1 U297 ( .A(n309), .Y(n173) );
  AND2X1 U299 ( .A(fifo_array[119]), .B(n5835), .Y(n303) );
  INVX1 U301 ( .A(n303), .Y(n174) );
  AND2X1 U303 ( .A(fifo_array[83]), .B(n5836), .Y(n265) );
  INVX1 U305 ( .A(n265), .Y(n175) );
  AND2X1 U307 ( .A(fifo_array[77]), .B(n5837), .Y(n259) );
  INVX1 U309 ( .A(n259), .Y(n176) );
  AND2X1 U311 ( .A(fifo_array[41]), .B(n5839), .Y(n220) );
  INVX1 U313 ( .A(n220), .Y(n177) );
  AND2X1 U315 ( .A(fifo_array[35]), .B(n5839), .Y(n214) );
  INVX1 U317 ( .A(n214), .Y(n1585) );
  AND2X1 U319 ( .A(fifo_array[1341]), .B(n5777), .Y(n1563) );
  INVX1 U321 ( .A(n1563), .Y(n3013) );
  AND2X1 U323 ( .A(fifo_array[1325]), .B(n5776), .Y(n1547) );
  INVX1 U325 ( .A(n1547), .Y(n3014) );
  AND2X1 U327 ( .A(fifo_array[1313]), .B(n5776), .Y(n1535) );
  INVX1 U329 ( .A(n1535), .Y(n3015) );
  AND2X1 U331 ( .A(fifo_array[1290]), .B(n5778), .Y(n1511) );
  INVX1 U333 ( .A(n1511), .Y(n3016) );
  AND2X1 U335 ( .A(fifo_array[1284]), .B(n5778), .Y(n1505) );
  INVX1 U337 ( .A(n1505), .Y(n3017) );
  AND2X1 U339 ( .A(fifo_array[1272]), .B(n5779), .Y(n1493) );
  INVX1 U341 ( .A(n1493), .Y(n3018) );
  AND2X1 U343 ( .A(fifo_array[1255]), .B(n5781), .Y(n1475) );
  INVX1 U345 ( .A(n1475), .Y(n3019) );
  AND2X1 U347 ( .A(fifo_array[1249]), .B(n5780), .Y(n1469) );
  INVX1 U349 ( .A(n1469), .Y(n3020) );
  AND2X1 U351 ( .A(fifo_array[1214]), .B(n5783), .Y(n1433) );
  INVX1 U353 ( .A(n1433), .Y(n3021) );
  AND2X1 U355 ( .A(fifo_array[1208]), .B(n5782), .Y(n1427) );
  INVX1 U357 ( .A(n1427), .Y(n3022) );
  AND2X1 U359 ( .A(fifo_array[1167]), .B(n5784), .Y(n1385) );
  INVX1 U361 ( .A(n1385), .Y(n3023) );
  AND2X1 U363 ( .A(fifo_array[1132]), .B(n5787), .Y(n1349) );
  INVX1 U365 ( .A(n1349), .Y(n3024) );
  AND2X1 U367 ( .A(fifo_array[1126]), .B(n5786), .Y(n1343) );
  INVX1 U369 ( .A(n1343), .Y(n3025) );
  AND2X1 U371 ( .A(fifo_array[1065]), .B(n5788), .Y(n1281) );
  INVX1 U372 ( .A(n1281), .Y(n3026) );
  AND2X1 U374 ( .A(fifo_array[1053]), .B(n5789), .Y(n1269) );
  INVX1 U376 ( .A(n1269), .Y(n3027) );
  AND2X1 U378 ( .A(fifo_array[1025]), .B(n5790), .Y(n1239) );
  INVX1 U380 ( .A(n1239), .Y(n3028) );
  AND2X1 U382 ( .A(fifo_array[1012]), .B(n5791), .Y(n1226) );
  INVX1 U384 ( .A(n1226), .Y(n3029) );
  AND2X1 U386 ( .A(fifo_array[993]), .B(n5793), .Y(n1206) );
  INVX1 U388 ( .A(n1206), .Y(n3030) );
  AND2X1 U390 ( .A(fifo_array[984]), .B(n5792), .Y(n1197) );
  INVX1 U392 ( .A(n1197), .Y(n3031) );
  AND2X1 U394 ( .A(fifo_array[971]), .B(n5792), .Y(n1184) );
  INVX1 U396 ( .A(n1184), .Y(n3032) );
  AND2X1 U398 ( .A(fifo_array[952]), .B(n5795), .Y(n1164) );
  INVX1 U400 ( .A(n1164), .Y(n3033) );
  AND2X1 U402 ( .A(fifo_array[943]), .B(n5794), .Y(n1155) );
  INVX1 U404 ( .A(n1155), .Y(n3034) );
  AND2X1 U406 ( .A(fifo_array[930]), .B(n5794), .Y(n1142) );
  INVX1 U408 ( .A(n1142), .Y(n3035) );
  AND2X1 U410 ( .A(fifo_array[911]), .B(n5797), .Y(n1122) );
  INVX1 U412 ( .A(n1122), .Y(n3036) );
  AND2X1 U414 ( .A(fifo_array[902]), .B(n5796), .Y(n1113) );
  INVX1 U416 ( .A(n1113), .Y(n3037) );
  AND2X1 U418 ( .A(fifo_array[889]), .B(n5796), .Y(n1100) );
  INVX1 U420 ( .A(n1100), .Y(n3038) );
  AND2X1 U422 ( .A(fifo_array[856]), .B(n5799), .Y(n1066) );
  INVX1 U424 ( .A(n1066), .Y(n3039) );
  AND2X1 U426 ( .A(fifo_array[849]), .B(n5799), .Y(n1059) );
  INVX1 U428 ( .A(n1059), .Y(n3040) );
  AND2X1 U430 ( .A(fifo_array[834]), .B(n5801), .Y(n1043) );
  INVX1 U432 ( .A(n1043), .Y(n3041) );
  AND2X1 U434 ( .A(fifo_array[820]), .B(n5800), .Y(n1029) );
  INVX1 U436 ( .A(n1029), .Y(n3042) );
  AND2X1 U438 ( .A(fifo_array[808]), .B(n5801), .Y(n1017) );
  INVX1 U440 ( .A(n1017), .Y(n3043) );
  AND2X1 U442 ( .A(fifo_array[795]), .B(n5803), .Y(n1003) );
  INVX1 U444 ( .A(n1003), .Y(n3044) );
  AND2X1 U446 ( .A(fifo_array[779]), .B(n5802), .Y(n987) );
  INVX1 U448 ( .A(n987), .Y(n3045) );
  AND2X1 U450 ( .A(fifo_array[767]), .B(n5803), .Y(n975) );
  INVX1 U452 ( .A(n975), .Y(n3046) );
  AND2X1 U454 ( .A(fifo_array[744]), .B(n5805), .Y(n951) );
  INVX1 U456 ( .A(n951), .Y(n3047) );
  AND2X1 U457 ( .A(fifo_array[738]), .B(n5804), .Y(n945) );
  INVX1 U459 ( .A(n945), .Y(n3048) );
  AND2X1 U461 ( .A(fifo_array[726]), .B(n5804), .Y(n933) );
  INVX1 U463 ( .A(n933), .Y(n3049) );
  AND2X1 U465 ( .A(fifo_array[709]), .B(n5807), .Y(n914) );
  INVX1 U467 ( .A(n914), .Y(n3050) );
  AND2X1 U469 ( .A(fifo_array[703]), .B(n5807), .Y(n908) );
  INVX1 U471 ( .A(n908), .Y(n3051) );
  AND2X1 U473 ( .A(fifo_array[668]), .B(n5809), .Y(n872) );
  INVX1 U475 ( .A(n872), .Y(n3052) );
  AND2X1 U477 ( .A(fifo_array[662]), .B(n5809), .Y(n866) );
  INVX1 U479 ( .A(n866), .Y(n3053) );
  AND2X1 U481 ( .A(fifo_array[621]), .B(n5811), .Y(n824) );
  INVX1 U483 ( .A(n824), .Y(n3054) );
  AND2X1 U485 ( .A(fifo_array[586]), .B(n5813), .Y(n788) );
  INVX1 U487 ( .A(n788), .Y(n3055) );
  AND2X1 U489 ( .A(fifo_array[580]), .B(n5813), .Y(n782) );
  INVX1 U491 ( .A(n782), .Y(n3056) );
  AND2X1 U493 ( .A(fifo_array[519]), .B(n5815), .Y(n720) );
  INVX1 U495 ( .A(n720), .Y(n3057) );
  AND2X1 U497 ( .A(fifo_array[507]), .B(n5814), .Y(n708) );
  INVX1 U499 ( .A(n708), .Y(n3058) );
  AND2X1 U501 ( .A(fifo_array[479]), .B(n5817), .Y(n679) );
  INVX1 U503 ( .A(n679), .Y(n3059) );
  AND2X1 U505 ( .A(fifo_array[466]), .B(n5816), .Y(n666) );
  INVX1 U507 ( .A(n666), .Y(n3060) );
  AND2X1 U509 ( .A(fifo_array[447]), .B(n5819), .Y(n646) );
  INVX1 U511 ( .A(n646), .Y(n3061) );
  AND2X1 U513 ( .A(fifo_array[438]), .B(n5818), .Y(n637) );
  INVX1 U515 ( .A(n637), .Y(n3062) );
  AND2X1 U517 ( .A(fifo_array[425]), .B(n5818), .Y(n624) );
  INVX1 U519 ( .A(n624), .Y(n3063) );
  AND2X1 U521 ( .A(fifo_array[406]), .B(n5821), .Y(n604) );
  INVX1 U523 ( .A(n604), .Y(n3064) );
  AND2X1 U525 ( .A(fifo_array[397]), .B(n5820), .Y(n595) );
  INVX1 U527 ( .A(n595), .Y(n3065) );
  AND2X1 U529 ( .A(fifo_array[384]), .B(n5820), .Y(n582) );
  INVX1 U531 ( .A(n582), .Y(n3066) );
  AND2X1 U533 ( .A(fifo_array[365]), .B(n5823), .Y(n561) );
  INVX1 U535 ( .A(n561), .Y(n3067) );
  AND2X1 U537 ( .A(fifo_array[356]), .B(n5822), .Y(n552) );
  INVX1 U539 ( .A(n552), .Y(n3068) );
  AND2X1 U541 ( .A(fifo_array[343]), .B(n5822), .Y(n539) );
  INVX1 U542 ( .A(n539), .Y(n3069) );
  AND2X1 U544 ( .A(fifo_array[310]), .B(n5825), .Y(n504) );
  INVX1 U546 ( .A(n504), .Y(n3070) );
  AND2X1 U548 ( .A(fifo_array[303]), .B(n5825), .Y(n497) );
  INVX1 U550 ( .A(n497), .Y(n3071) );
  AND2X1 U552 ( .A(fifo_array[288]), .B(n5827), .Y(n480) );
  INVX1 U554 ( .A(n480), .Y(n3072) );
  AND2X1 U556 ( .A(fifo_array[274]), .B(n5826), .Y(n466) );
  INVX1 U558 ( .A(n466), .Y(n3073) );
  AND2X1 U560 ( .A(fifo_array[262]), .B(n5827), .Y(n454) );
  INVX1 U562 ( .A(n454), .Y(n3074) );
  AND2X1 U564 ( .A(fifo_array[249]), .B(n5829), .Y(n439) );
  INVX1 U566 ( .A(n439), .Y(n3075) );
  AND2X1 U568 ( .A(fifo_array[233]), .B(n5828), .Y(n423) );
  INVX1 U570 ( .A(n423), .Y(n3076) );
  AND2X1 U572 ( .A(fifo_array[221]), .B(n5829), .Y(n411) );
  INVX1 U574 ( .A(n411), .Y(n3077) );
  AND2X1 U576 ( .A(fifo_array[198]), .B(n5831), .Y(n386) );
  INVX1 U578 ( .A(n386), .Y(n3078) );
  AND2X1 U580 ( .A(fifo_array[192]), .B(n5830), .Y(n380) );
  INVX1 U582 ( .A(n380), .Y(n3079) );
  AND2X1 U584 ( .A(fifo_array[180]), .B(n5830), .Y(n368) );
  INVX1 U586 ( .A(n368), .Y(n3080) );
  AND2X1 U588 ( .A(fifo_array[163]), .B(n5833), .Y(n349) );
  INVX1 U590 ( .A(n349), .Y(n3081) );
  AND2X1 U592 ( .A(fifo_array[157]), .B(n5833), .Y(n343) );
  INVX1 U594 ( .A(n343), .Y(n3082) );
  AND2X1 U596 ( .A(fifo_array[122]), .B(n5835), .Y(n306) );
  INVX1 U598 ( .A(n306), .Y(n3083) );
  AND2X1 U600 ( .A(fifo_array[116]), .B(n5835), .Y(n300) );
  INVX1 U602 ( .A(n300), .Y(n3084) );
  AND2X1 U604 ( .A(fifo_array[75]), .B(n5837), .Y(n257) );
  INVX1 U606 ( .A(n257), .Y(n3085) );
  AND2X1 U608 ( .A(fifo_array[40]), .B(n5839), .Y(n219) );
  INVX1 U610 ( .A(n219), .Y(n3086) );
  AND2X1 U612 ( .A(fifo_array[34]), .B(n5838), .Y(n213) );
  INVX1 U614 ( .A(n213), .Y(n3087) );
  AND2X1 U616 ( .A(fifo_array[1332]), .B(n5776), .Y(n1554) );
  INVX1 U618 ( .A(n1554), .Y(n3088) );
  AND2X1 U620 ( .A(fifo_array[1326]), .B(n5777), .Y(n1548) );
  INVX1 U622 ( .A(n1548), .Y(n3089) );
  AND2X1 U624 ( .A(fifo_array[1314]), .B(n5777), .Y(n1536) );
  INVX1 U626 ( .A(n1536), .Y(n3090) );
  AND2X1 U627 ( .A(fifo_array[1299]), .B(n5779), .Y(n1520) );
  INVX1 U629 ( .A(n1520), .Y(n3091) );
  AND2X1 U631 ( .A(fifo_array[1283]), .B(n5779), .Y(n1504) );
  INVX1 U633 ( .A(n1504), .Y(n3092) );
  AND2X1 U635 ( .A(fifo_array[1271]), .B(n5778), .Y(n1492) );
  INVX1 U637 ( .A(n1492), .Y(n3093) );
  AND2X1 U639 ( .A(fifo_array[1256]), .B(n5781), .Y(n1476) );
  INVX1 U641 ( .A(n1476), .Y(n3094) );
  AND2X1 U643 ( .A(fifo_array[1250]), .B(n5780), .Y(n1470) );
  INVX1 U645 ( .A(n1470), .Y(n3095) );
  AND2X1 U647 ( .A(fifo_array[1213]), .B(n5783), .Y(n1432) );
  INVX1 U649 ( .A(n1432), .Y(n3096) );
  AND2X1 U651 ( .A(fifo_array[1207]), .B(n5782), .Y(n1426) );
  INVX1 U653 ( .A(n1426), .Y(n3097) );
  AND2X1 U655 ( .A(fifo_array[1174]), .B(n5785), .Y(n1392) );
  INVX1 U657 ( .A(n1392), .Y(n3098) );
  AND2X1 U659 ( .A(fifo_array[1168]), .B(n5784), .Y(n1386) );
  INVX1 U661 ( .A(n1386), .Y(n3099) );
  AND2X1 U663 ( .A(fifo_array[1125]), .B(n5786), .Y(n1342) );
  INVX1 U665 ( .A(n1342), .Y(n3100) );
  AND2X1 U667 ( .A(fifo_array[1076]), .B(n5789), .Y(n1292) );
  INVX1 U669 ( .A(n1292), .Y(n3101) );
  AND2X1 U671 ( .A(fifo_array[1064]), .B(n5789), .Y(n1280) );
  INVX1 U673 ( .A(n1280), .Y(n3102) );
  AND2X1 U675 ( .A(fifo_array[1052]), .B(n5789), .Y(n1268) );
  INVX1 U677 ( .A(n1268), .Y(n3103) );
  AND2X1 U679 ( .A(fifo_array[1035]), .B(n5791), .Y(n1249) );
  INVX1 U681 ( .A(n1249), .Y(n3104) );
  AND2X1 U683 ( .A(fifo_array[1026]), .B(n5791), .Y(n1240) );
  INVX1 U685 ( .A(n1240), .Y(n3105) );
  AND2X1 U687 ( .A(fifo_array[1013]), .B(n5791), .Y(n1227) );
  INVX1 U689 ( .A(n1227), .Y(n3106) );
  AND2X1 U691 ( .A(fifo_array[983]), .B(n5793), .Y(n1196) );
  INVX1 U693 ( .A(n1196), .Y(n3107) );
  AND2X1 U695 ( .A(fifo_array[970]), .B(n5792), .Y(n1183) );
  INVX1 U697 ( .A(n1183), .Y(n3108) );
  AND2X1 U699 ( .A(fifo_array[953]), .B(n5795), .Y(n1165) );
  INVX1 U701 ( .A(n1165), .Y(n3109) );
  AND2X1 U703 ( .A(fifo_array[944]), .B(n5794), .Y(n1156) );
  INVX1 U705 ( .A(n1156), .Y(n3110) );
  AND2X1 U707 ( .A(fifo_array[931]), .B(n5794), .Y(n1143) );
  INVX1 U709 ( .A(n1143), .Y(n3111) );
  AND2X1 U711 ( .A(fifo_array[910]), .B(n5797), .Y(n1121) );
  INVX1 U712 ( .A(n1121), .Y(n3112) );
  AND2X1 U714 ( .A(fifo_array[901]), .B(n5796), .Y(n1112) );
  INVX1 U716 ( .A(n1112), .Y(n3113) );
  AND2X1 U718 ( .A(fifo_array[888]), .B(n5796), .Y(n1099) );
  INVX1 U720 ( .A(n1099), .Y(n3114) );
  AND2X1 U722 ( .A(fifo_array[876]), .B(n5798), .Y(n1086) );
  INVX1 U724 ( .A(n1086), .Y(n3115) );
  AND2X1 U726 ( .A(fifo_array[862]), .B(n5798), .Y(n1072) );
  INVX1 U728 ( .A(n1072), .Y(n3116) );
  AND2X1 U730 ( .A(fifo_array[850]), .B(n5799), .Y(n1060) );
  INVX1 U732 ( .A(n1060), .Y(n3117) );
  AND2X1 U734 ( .A(fifo_array[814]), .B(n5800), .Y(n1023) );
  INVX1 U736 ( .A(n1023), .Y(n3118) );
  AND2X1 U738 ( .A(fifo_array[807]), .B(n5801), .Y(n1016) );
  INVX1 U740 ( .A(n1016), .Y(n3119) );
  AND2X1 U742 ( .A(fifo_array[786]), .B(n5803), .Y(n994) );
  INVX1 U744 ( .A(n994), .Y(n3120) );
  AND2X1 U746 ( .A(fifo_array[780]), .B(n5802), .Y(n988) );
  INVX1 U748 ( .A(n988), .Y(n3121) );
  AND2X1 U750 ( .A(fifo_array[768]), .B(n5802), .Y(n976) );
  INVX1 U752 ( .A(n976), .Y(n3122) );
  AND2X1 U754 ( .A(fifo_array[753]), .B(n5805), .Y(n960) );
  INVX1 U756 ( .A(n960), .Y(n3123) );
  AND2X1 U758 ( .A(fifo_array[737]), .B(n5804), .Y(n944) );
  INVX1 U760 ( .A(n944), .Y(n3124) );
  AND2X1 U762 ( .A(fifo_array[725]), .B(n5805), .Y(n932) );
  INVX1 U764 ( .A(n932), .Y(n3125) );
  AND2X1 U766 ( .A(fifo_array[710]), .B(n5806), .Y(n915) );
  INVX1 U768 ( .A(n915), .Y(n3126) );
  AND2X1 U770 ( .A(fifo_array[704]), .B(n5807), .Y(n909) );
  INVX1 U772 ( .A(n909), .Y(n3127) );
  AND2X1 U774 ( .A(fifo_array[667]), .B(n5808), .Y(n871) );
  INVX1 U776 ( .A(n871), .Y(n3128) );
  AND2X1 U778 ( .A(fifo_array[661]), .B(n5809), .Y(n865) );
  INVX1 U780 ( .A(n865), .Y(n3129) );
  AND2X1 U782 ( .A(fifo_array[628]), .B(n5811), .Y(n831) );
  INVX1 U784 ( .A(n831), .Y(n3130) );
  AND2X1 U786 ( .A(fifo_array[622]), .B(n5811), .Y(n825) );
  INVX1 U788 ( .A(n825), .Y(n3131) );
  AND2X1 U790 ( .A(fifo_array[579]), .B(n5813), .Y(n781) );
  INVX1 U792 ( .A(n781), .Y(n3132) );
  AND2X1 U794 ( .A(fifo_array[530]), .B(n5814), .Y(n731) );
  INVX1 U796 ( .A(n731), .Y(n3133) );
  AND2X1 U797 ( .A(fifo_array[518]), .B(n5815), .Y(n719) );
  INVX1 U800 ( .A(n719), .Y(n3134) );
  AND2X1 U802 ( .A(fifo_array[506]), .B(n5814), .Y(n707) );
  INVX1 U804 ( .A(n707), .Y(n3135) );
  AND2X1 U806 ( .A(fifo_array[489]), .B(n5817), .Y(n689) );
  INVX1 U808 ( .A(n689), .Y(n3136) );
  AND2X1 U810 ( .A(fifo_array[480]), .B(n5816), .Y(n680) );
  INVX1 U812 ( .A(n680), .Y(n3137) );
  AND2X1 U814 ( .A(fifo_array[467]), .B(n5816), .Y(n667) );
  INVX1 U816 ( .A(n667), .Y(n3138) );
  AND2X1 U818 ( .A(fifo_array[437]), .B(n5819), .Y(n636) );
  INVX1 U820 ( .A(n636), .Y(n3139) );
  AND2X1 U822 ( .A(fifo_array[424]), .B(n5818), .Y(n623) );
  INVX1 U824 ( .A(n623), .Y(n3140) );
  AND2X1 U826 ( .A(fifo_array[407]), .B(n5821), .Y(n605) );
  INVX1 U828 ( .A(n605), .Y(n3141) );
  AND2X1 U830 ( .A(fifo_array[398]), .B(n5820), .Y(n596) );
  INVX1 U832 ( .A(n596), .Y(n3142) );
  AND2X1 U834 ( .A(fifo_array[385]), .B(n5820), .Y(n583) );
  INVX1 U836 ( .A(n583), .Y(n3143) );
  AND2X1 U838 ( .A(fifo_array[364]), .B(n5823), .Y(n560) );
  INVX1 U840 ( .A(n560), .Y(n3144) );
  AND2X1 U842 ( .A(fifo_array[355]), .B(n5822), .Y(n551) );
  INVX1 U844 ( .A(n551), .Y(n3145) );
  AND2X1 U846 ( .A(fifo_array[342]), .B(n5822), .Y(n538) );
  INVX1 U848 ( .A(n538), .Y(n3146) );
  AND2X1 U850 ( .A(fifo_array[330]), .B(n5824), .Y(n524) );
  INVX1 U852 ( .A(n524), .Y(n3147) );
  AND2X1 U854 ( .A(fifo_array[316]), .B(n5824), .Y(n510) );
  INVX1 U856 ( .A(n510), .Y(n3148) );
  AND2X1 U858 ( .A(fifo_array[304]), .B(n5825), .Y(n498) );
  INVX1 U860 ( .A(n498), .Y(n3149) );
  AND2X1 U862 ( .A(fifo_array[268]), .B(n5826), .Y(n460) );
  INVX1 U864 ( .A(n460), .Y(n3150) );
  AND2X1 U866 ( .A(fifo_array[261]), .B(n5827), .Y(n453) );
  INVX1 U868 ( .A(n453), .Y(n3151) );
  AND2X1 U870 ( .A(fifo_array[240]), .B(n5829), .Y(n430) );
  INVX1 U872 ( .A(n430), .Y(n3152) );
  AND2X1 U874 ( .A(fifo_array[234]), .B(n5828), .Y(n424) );
  INVX1 U876 ( .A(n424), .Y(n3153) );
  AND2X1 U878 ( .A(fifo_array[222]), .B(n5828), .Y(n412) );
  INVX1 U880 ( .A(n412), .Y(n3154) );
  AND2X1 U882 ( .A(fifo_array[207]), .B(n5831), .Y(n395) );
  INVX1 U883 ( .A(n395), .Y(n3155) );
  AND2X1 U885 ( .A(fifo_array[191]), .B(n5830), .Y(n379) );
  INVX1 U887 ( .A(n379), .Y(n3156) );
  AND2X1 U889 ( .A(fifo_array[179]), .B(n5831), .Y(n367) );
  INVX1 U891 ( .A(n367), .Y(n3157) );
  AND2X1 U893 ( .A(fifo_array[164]), .B(n5832), .Y(n350) );
  INVX1 U895 ( .A(n350), .Y(n3158) );
  AND2X1 U897 ( .A(fifo_array[158]), .B(n5833), .Y(n344) );
  INVX1 U899 ( .A(n344), .Y(n3159) );
  AND2X1 U901 ( .A(fifo_array[121]), .B(n5834), .Y(n305) );
  INVX1 U903 ( .A(n305), .Y(n3160) );
  AND2X1 U905 ( .A(fifo_array[115]), .B(n5835), .Y(n299) );
  INVX1 U907 ( .A(n299), .Y(n3161) );
  AND2X1 U909 ( .A(fifo_array[82]), .B(n5837), .Y(n264) );
  INVX1 U911 ( .A(n264), .Y(n3162) );
  AND2X1 U913 ( .A(fifo_array[76]), .B(n5837), .Y(n258) );
  INVX1 U915 ( .A(n258), .Y(n3163) );
  AND2X1 U917 ( .A(fifo_array[33]), .B(n5838), .Y(n212) );
  INVX1 U919 ( .A(n212), .Y(n3164) );
  AND2X1 U921 ( .A(fifo_array[1318]), .B(n5777), .Y(n1540) );
  INVX1 U923 ( .A(n1540), .Y(n3165) );
  AND2X1 U925 ( .A(fifo_array[1311]), .B(n5776), .Y(n1533) );
  INVX1 U927 ( .A(n1533), .Y(n3166) );
  AND2X1 U929 ( .A(fifo_array[1296]), .B(n5779), .Y(n1517) );
  INVX1 U931 ( .A(n1517), .Y(n3167) );
  AND2X1 U933 ( .A(fifo_array[1282]), .B(n5778), .Y(n1503) );
  INVX1 U935 ( .A(n1503), .Y(n3168) );
  AND2X1 U937 ( .A(fifo_array[1270]), .B(n5778), .Y(n1491) );
  INVX1 U939 ( .A(n1491), .Y(n3169) );
  AND2X1 U941 ( .A(fifo_array[1251]), .B(n5780), .Y(n1471) );
  INVX1 U943 ( .A(n1471), .Y(n3170) );
  AND2X1 U945 ( .A(fifo_array[1216]), .B(n5783), .Y(n1435) );
  INVX1 U947 ( .A(n1435), .Y(n3171) );
  AND2X1 U949 ( .A(fifo_array[1210]), .B(n5782), .Y(n1429) );
  INVX1 U951 ( .A(n1429), .Y(n3172) );
  AND2X1 U953 ( .A(fifo_array[1171]), .B(n5785), .Y(n1389) );
  INVX1 U955 ( .A(n1389), .Y(n3173) );
  AND2X1 U957 ( .A(fifo_array[1165]), .B(n5784), .Y(n1383) );
  INVX1 U959 ( .A(n1383), .Y(n3174) );
  AND2X1 U961 ( .A(fifo_array[1130]), .B(n5787), .Y(n1347) );
  INVX1 U963 ( .A(n1347), .Y(n3175) );
  AND2X1 U965 ( .A(fifo_array[1124]), .B(n5786), .Y(n1341) );
  INVX1 U967 ( .A(n1341), .Y(n3176) );
  AND2X1 U968 ( .A(fifo_array[1075]), .B(n5788), .Y(n1291) );
  INVX1 U970 ( .A(n1291), .Y(n3177) );
  AND2X1 U972 ( .A(fifo_array[1063]), .B(n5789), .Y(n1279) );
  INVX1 U974 ( .A(n1279), .Y(n3178) );
  AND2X1 U976 ( .A(fifo_array[1051]), .B(n5789), .Y(n1267) );
  INVX1 U978 ( .A(n1267), .Y(n3179) );
  AND2X1 U980 ( .A(fifo_array[1036]), .B(n5790), .Y(n1250) );
  INVX1 U982 ( .A(n1250), .Y(n3180) );
  AND2X1 U984 ( .A(fifo_array[1027]), .B(n5790), .Y(n1241) );
  INVX1 U986 ( .A(n1241), .Y(n3181) );
  AND2X1 U988 ( .A(fifo_array[1014]), .B(n5791), .Y(n1228) );
  INVX1 U990 ( .A(n1228), .Y(n3182) );
  AND2X1 U992 ( .A(fifo_array[995]), .B(n5793), .Y(n1208) );
  INVX1 U994 ( .A(n1208), .Y(n3183) );
  AND2X1 U996 ( .A(fifo_array[986]), .B(n5792), .Y(n1199) );
  INVX1 U998 ( .A(n1199), .Y(n3184) );
  AND2X1 U1000 ( .A(fifo_array[973]), .B(n5792), .Y(n1186) );
  INVX1 U1002 ( .A(n1186), .Y(n3185) );
  AND2X1 U1004 ( .A(fifo_array[941]), .B(n5795), .Y(n1153) );
  INVX1 U1006 ( .A(n1153), .Y(n3186) );
  AND2X1 U1008 ( .A(fifo_array[928]), .B(n5794), .Y(n1140) );
  INVX1 U1010 ( .A(n1140), .Y(n3187) );
  AND2X1 U1012 ( .A(fifo_array[909]), .B(n5797), .Y(n1120) );
  INVX1 U1014 ( .A(n1120), .Y(n3188) );
  AND2X1 U1016 ( .A(fifo_array[900]), .B(n5796), .Y(n1111) );
  INVX1 U1018 ( .A(n1111), .Y(n3189) );
  AND2X1 U1020 ( .A(fifo_array[887]), .B(n5796), .Y(n1098) );
  INVX1 U1022 ( .A(n1098), .Y(n3190) );
  AND2X1 U1024 ( .A(fifo_array[879]), .B(n5799), .Y(n1089) );
  INVX1 U1026 ( .A(n1089), .Y(n3191) );
  AND2X1 U1028 ( .A(fifo_array[863]), .B(n5798), .Y(n1073) );
  INVX1 U1030 ( .A(n1073), .Y(n3192) );
  AND2X1 U1032 ( .A(fifo_array[851]), .B(n5799), .Y(n1061) );
  INVX1 U1034 ( .A(n1061), .Y(n3193) );
  AND2X1 U1036 ( .A(fifo_array[828]), .B(n5801), .Y(n1037) );
  INVX1 U1038 ( .A(n1037), .Y(n3194) );
  AND2X1 U1040 ( .A(fifo_array[822]), .B(n5800), .Y(n1031) );
  INVX1 U1042 ( .A(n1031), .Y(n3195) );
  AND2X1 U1044 ( .A(fifo_array[810]), .B(n5800), .Y(n1019) );
  INVX1 U1046 ( .A(n1019), .Y(n3196) );
  AND2X1 U1048 ( .A(fifo_array[772]), .B(n5802), .Y(n980) );
  INVX1 U1050 ( .A(n980), .Y(n3197) );
  AND2X1 U1052 ( .A(fifo_array[765]), .B(n5803), .Y(n973) );
  INVX1 U1053 ( .A(n973), .Y(n3198) );
  AND2X1 U1055 ( .A(fifo_array[750]), .B(n5804), .Y(n957) );
  INVX1 U1057 ( .A(n957), .Y(n3199) );
  AND2X1 U1059 ( .A(fifo_array[736]), .B(n5804), .Y(n943) );
  INVX1 U1061 ( .A(n943), .Y(n3200) );
  AND2X1 U1063 ( .A(fifo_array[724]), .B(n5805), .Y(n931) );
  INVX1 U1065 ( .A(n931), .Y(n3201) );
  AND2X1 U1067 ( .A(fifo_array[705]), .B(n5807), .Y(n910) );
  INVX1 U1069 ( .A(n910), .Y(n3202) );
  AND2X1 U1071 ( .A(fifo_array[670]), .B(n5809), .Y(n874) );
  INVX1 U1073 ( .A(n874), .Y(n3203) );
  AND2X1 U1075 ( .A(fifo_array[664]), .B(n5809), .Y(n868) );
  INVX1 U1077 ( .A(n868), .Y(n3204) );
  AND2X1 U1079 ( .A(fifo_array[625]), .B(n5810), .Y(n828) );
  INVX1 U1081 ( .A(n828), .Y(n3205) );
  AND2X1 U1083 ( .A(fifo_array[619]), .B(n5811), .Y(n822) );
  INVX1 U1085 ( .A(n822), .Y(n3206) );
  AND2X1 U1087 ( .A(fifo_array[584]), .B(n5812), .Y(n786) );
  INVX1 U1089 ( .A(n786), .Y(n3207) );
  AND2X1 U1091 ( .A(fifo_array[578]), .B(n5813), .Y(n780) );
  INVX1 U1093 ( .A(n780), .Y(n3208) );
  AND2X1 U1095 ( .A(fifo_array[529]), .B(n5814), .Y(n730) );
  INVX1 U1097 ( .A(n730), .Y(n3209) );
  AND2X1 U1099 ( .A(fifo_array[517]), .B(n5815), .Y(n718) );
  INVX1 U1101 ( .A(n718), .Y(n3210) );
  AND2X1 U1103 ( .A(fifo_array[505]), .B(n5815), .Y(n706) );
  INVX1 U1105 ( .A(n706), .Y(n3211) );
  AND2X1 U1107 ( .A(fifo_array[490]), .B(n5817), .Y(n690) );
  INVX1 U1109 ( .A(n690), .Y(n3212) );
  AND2X1 U1111 ( .A(fifo_array[481]), .B(n5816), .Y(n681) );
  INVX1 U1113 ( .A(n681), .Y(n3213) );
  AND2X1 U1115 ( .A(fifo_array[468]), .B(n5816), .Y(n668) );
  INVX1 U1117 ( .A(n668), .Y(n3214) );
  AND2X1 U1119 ( .A(fifo_array[449]), .B(n5819), .Y(n648) );
  INVX1 U1121 ( .A(n648), .Y(n3215) );
  AND2X1 U1123 ( .A(fifo_array[440]), .B(n5818), .Y(n639) );
  INVX1 U1125 ( .A(n639), .Y(n3216) );
  AND2X1 U1127 ( .A(fifo_array[427]), .B(n5818), .Y(n626) );
  INVX1 U1129 ( .A(n626), .Y(n3217) );
  AND2X1 U1131 ( .A(fifo_array[395]), .B(n5821), .Y(n593) );
  INVX1 U1133 ( .A(n593), .Y(n3218) );
  AND2X1 U1135 ( .A(fifo_array[382]), .B(n5820), .Y(n580) );
  INVX1 U1137 ( .A(n580), .Y(n3219) );
  AND2X1 U1138 ( .A(fifo_array[363]), .B(n5823), .Y(n559) );
  INVX1 U1140 ( .A(n559), .Y(n3220) );
  AND2X1 U1142 ( .A(fifo_array[354]), .B(n5822), .Y(n550) );
  INVX1 U1144 ( .A(n550), .Y(n3221) );
  AND2X1 U1146 ( .A(fifo_array[341]), .B(n5822), .Y(n537) );
  INVX1 U1148 ( .A(n537), .Y(n3222) );
  AND2X1 U1150 ( .A(fifo_array[333]), .B(n5825), .Y(n527) );
  INVX1 U1152 ( .A(n527), .Y(n3223) );
  AND2X1 U1154 ( .A(fifo_array[317]), .B(n5824), .Y(n511) );
  INVX1 U1156 ( .A(n511), .Y(n3224) );
  AND2X1 U1158 ( .A(fifo_array[305]), .B(n5825), .Y(n499) );
  INVX1 U1160 ( .A(n499), .Y(n3225) );
  AND2X1 U1162 ( .A(fifo_array[282]), .B(n5827), .Y(n474) );
  INVX1 U1164 ( .A(n474), .Y(n3226) );
  AND2X1 U1166 ( .A(fifo_array[276]), .B(n5826), .Y(n468) );
  INVX1 U1168 ( .A(n468), .Y(n3227) );
  AND2X1 U1170 ( .A(fifo_array[264]), .B(n5826), .Y(n456) );
  INVX1 U1172 ( .A(n456), .Y(n3228) );
  AND2X1 U1174 ( .A(fifo_array[226]), .B(n5828), .Y(n416) );
  INVX1 U1176 ( .A(n416), .Y(n3229) );
  AND2X1 U1178 ( .A(fifo_array[219]), .B(n5829), .Y(n409) );
  INVX1 U1180 ( .A(n409), .Y(n3230) );
  AND2X1 U1182 ( .A(fifo_array[204]), .B(n5830), .Y(n392) );
  INVX1 U1184 ( .A(n392), .Y(n3231) );
  AND2X1 U1186 ( .A(fifo_array[190]), .B(n5830), .Y(n378) );
  INVX1 U1188 ( .A(n378), .Y(n3232) );
  AND2X1 U1190 ( .A(fifo_array[178]), .B(n5831), .Y(n366) );
  INVX1 U1192 ( .A(n366), .Y(n3233) );
  AND2X1 U1194 ( .A(fifo_array[159]), .B(n5833), .Y(n345) );
  INVX1 U1196 ( .A(n345), .Y(n3234) );
  AND2X1 U1198 ( .A(fifo_array[124]), .B(n5835), .Y(n308) );
  INVX1 U1200 ( .A(n308), .Y(n3235) );
  AND2X1 U1202 ( .A(fifo_array[118]), .B(n5835), .Y(n302) );
  INVX1 U1204 ( .A(n302), .Y(n3236) );
  AND2X1 U1206 ( .A(fifo_array[79]), .B(n5836), .Y(n261) );
  INVX1 U1208 ( .A(n261), .Y(n3237) );
  AND2X1 U1210 ( .A(fifo_array[73]), .B(n5837), .Y(n255) );
  INVX1 U1212 ( .A(n255), .Y(n3238) );
  AND2X1 U1214 ( .A(fifo_array[38]), .B(n5839), .Y(n217) );
  INVX1 U1216 ( .A(n217), .Y(n3239) );
  AND2X1 U1218 ( .A(fifo_array[32]), .B(n5839), .Y(n211) );
  INVX1 U1220 ( .A(n211), .Y(n3240) );
  AND2X1 U1222 ( .A(fifo_array[1338]), .B(n5777), .Y(n1560) );
  INVX1 U1223 ( .A(n1560), .Y(n3241) );
  AND2X1 U1225 ( .A(fifo_array[1324]), .B(n5776), .Y(n1546) );
  INVX1 U1227 ( .A(n1546), .Y(n3242) );
  AND2X1 U1229 ( .A(fifo_array[1312]), .B(n5776), .Y(n1534) );
  INVX1 U1231 ( .A(n1534), .Y(n3243) );
  AND2X1 U1233 ( .A(fifo_array[1276]), .B(n5779), .Y(n1497) );
  INVX1 U1235 ( .A(n1497), .Y(n3244) );
  AND2X1 U1237 ( .A(fifo_array[1269]), .B(n5778), .Y(n1490) );
  INVX1 U1239 ( .A(n1490), .Y(n3245) );
  AND2X1 U1241 ( .A(fifo_array[1258]), .B(n5781), .Y(n1478) );
  INVX1 U1243 ( .A(n1478), .Y(n3246) );
  AND2X1 U1245 ( .A(fifo_array[1252]), .B(n5780), .Y(n1472) );
  INVX1 U1247 ( .A(n1472), .Y(n3247) );
  AND2X1 U1249 ( .A(fifo_array[1209]), .B(n5782), .Y(n1428) );
  INVX1 U1251 ( .A(n1428), .Y(n3248) );
  AND2X1 U1253 ( .A(fifo_array[1172]), .B(n5785), .Y(n1390) );
  INVX1 U1255 ( .A(n1390), .Y(n3249) );
  AND2X1 U1257 ( .A(fifo_array[1166]), .B(n5784), .Y(n1384) );
  INVX1 U1259 ( .A(n1384), .Y(n3250) );
  AND2X1 U1261 ( .A(fifo_array[1129]), .B(n5787), .Y(n1346) );
  INVX1 U1263 ( .A(n1346), .Y(n3251) );
  AND2X1 U1265 ( .A(fifo_array[1123]), .B(n5786), .Y(n1340) );
  INVX1 U1267 ( .A(n1340), .Y(n3252) );
  AND2X1 U1269 ( .A(fifo_array[1071]), .B(n5789), .Y(n1287) );
  INVX1 U1271 ( .A(n1287), .Y(n3253) );
  AND2X1 U1273 ( .A(fifo_array[1058]), .B(n5788), .Y(n1274) );
  INVX1 U1275 ( .A(n1274), .Y(n3254) );
  AND2X1 U1277 ( .A(fifo_array[1050]), .B(n5789), .Y(n1266) );
  INVX1 U1279 ( .A(n1266), .Y(n3255) );
  AND2X1 U1281 ( .A(fifo_array[1037]), .B(n5791), .Y(n1251) );
  INVX1 U1283 ( .A(n1251), .Y(n3256) );
  AND2X1 U1285 ( .A(fifo_array[1028]), .B(n5791), .Y(n1242) );
  INVX1 U1287 ( .A(n1242), .Y(n3257) );
  AND2X1 U1289 ( .A(fifo_array[1015]), .B(n5791), .Y(n1229) );
  INVX1 U1291 ( .A(n1229), .Y(n3258) );
  AND2X1 U1293 ( .A(fifo_array[994]), .B(n5793), .Y(n1207) );
  INVX1 U1295 ( .A(n1207), .Y(n3259) );
  AND2X1 U1297 ( .A(fifo_array[985]), .B(n5792), .Y(n1198) );
  INVX1 U1299 ( .A(n1198), .Y(n3260) );
  AND2X1 U1301 ( .A(fifo_array[972]), .B(n5792), .Y(n1185) );
  INVX1 U1303 ( .A(n1185), .Y(n3261) );
  AND2X1 U1305 ( .A(fifo_array[951]), .B(n5795), .Y(n1163) );
  INVX1 U1307 ( .A(n1163), .Y(n3262) );
  AND2X1 U1308 ( .A(fifo_array[942]), .B(n5794), .Y(n1154) );
  INVX1 U1310 ( .A(n1154), .Y(n3263) );
  AND2X1 U1312 ( .A(fifo_array[929]), .B(n5794), .Y(n1141) );
  INVX1 U1314 ( .A(n1141), .Y(n3264) );
  AND2X1 U1316 ( .A(fifo_array[899]), .B(n5797), .Y(n1110) );
  INVX1 U1318 ( .A(n1110), .Y(n3265) );
  AND2X1 U1320 ( .A(fifo_array[886]), .B(n5796), .Y(n1097) );
  INVX1 U1322 ( .A(n1097), .Y(n3266) );
  AND2X1 U1324 ( .A(fifo_array[870]), .B(n5799), .Y(n1080) );
  INVX1 U1326 ( .A(n1080), .Y(n3267) );
  AND2X1 U1328 ( .A(fifo_array[864]), .B(n5798), .Y(n1074) );
  INVX1 U1330 ( .A(n1074), .Y(n3268) );
  AND2X1 U1332 ( .A(fifo_array[852]), .B(n5798), .Y(n1062) );
  INVX1 U1334 ( .A(n1062), .Y(n3269) );
  AND2X1 U1336 ( .A(fifo_array[837]), .B(n5801), .Y(n1046) );
  INVX1 U1338 ( .A(n1046), .Y(n3270) );
  AND2X1 U1340 ( .A(fifo_array[821]), .B(n5800), .Y(n1030) );
  INVX1 U1342 ( .A(n1030), .Y(n3271) );
  AND2X1 U1344 ( .A(fifo_array[809]), .B(n5801), .Y(n1018) );
  INVX1 U1346 ( .A(n1018), .Y(n3272) );
  AND2X1 U1348 ( .A(fifo_array[792]), .B(n5803), .Y(n1000) );
  INVX1 U1350 ( .A(n1000), .Y(n3273) );
  AND2X1 U1352 ( .A(fifo_array[778]), .B(n5802), .Y(n986) );
  INVX1 U1354 ( .A(n986), .Y(n3274) );
  AND2X1 U1356 ( .A(fifo_array[766]), .B(n5803), .Y(n974) );
  INVX1 U1358 ( .A(n974), .Y(n3275) );
  AND2X1 U1360 ( .A(fifo_array[730]), .B(n5805), .Y(n937) );
  INVX1 U1362 ( .A(n937), .Y(n3276) );
  AND2X1 U1364 ( .A(fifo_array[723]), .B(n5805), .Y(n930) );
  INVX1 U1366 ( .A(n930), .Y(n3277) );
  AND2X1 U1368 ( .A(fifo_array[712]), .B(n5807), .Y(n917) );
  INVX1 U1370 ( .A(n917), .Y(n3278) );
  AND2X1 U1372 ( .A(fifo_array[706]), .B(n5807), .Y(n911) );
  INVX1 U1374 ( .A(n911), .Y(n3279) );
  AND2X1 U1376 ( .A(fifo_array[663]), .B(n5809), .Y(n867) );
  INVX1 U1378 ( .A(n867), .Y(n3280) );
  AND2X1 U1380 ( .A(fifo_array[626]), .B(n5811), .Y(n829) );
  INVX1 U1382 ( .A(n829), .Y(n3281) );
  AND2X1 U1384 ( .A(fifo_array[620]), .B(n5811), .Y(n823) );
  INVX1 U1386 ( .A(n823), .Y(n3282) );
  AND2X1 U1388 ( .A(fifo_array[583]), .B(n5813), .Y(n785) );
  INVX1 U1390 ( .A(n785), .Y(n3283) );
  AND2X1 U1392 ( .A(fifo_array[577]), .B(n5813), .Y(n779) );
  INVX1 U1393 ( .A(n779), .Y(n3284) );
  AND2X1 U1395 ( .A(fifo_array[525]), .B(n5814), .Y(n726) );
  INVX1 U1397 ( .A(n726), .Y(n3285) );
  AND2X1 U1399 ( .A(fifo_array[512]), .B(n5815), .Y(n713) );
  INVX1 U1401 ( .A(n713), .Y(n3286) );
  AND2X1 U1403 ( .A(fifo_array[504]), .B(n5815), .Y(n705) );
  INVX1 U1405 ( .A(n705), .Y(n3287) );
  AND2X1 U1407 ( .A(fifo_array[491]), .B(n5817), .Y(n691) );
  INVX1 U1409 ( .A(n691), .Y(n3288) );
  AND2X1 U1411 ( .A(fifo_array[482]), .B(n5816), .Y(n682) );
  INVX1 U1413 ( .A(n682), .Y(n3289) );
  AND2X1 U1415 ( .A(fifo_array[469]), .B(n5816), .Y(n669) );
  INVX1 U1417 ( .A(n669), .Y(n3290) );
  AND2X1 U1419 ( .A(fifo_array[448]), .B(n5819), .Y(n647) );
  INVX1 U1421 ( .A(n647), .Y(n3291) );
  AND2X1 U1423 ( .A(fifo_array[439]), .B(n5818), .Y(n638) );
  INVX1 U1425 ( .A(n638), .Y(n3292) );
  AND2X1 U1427 ( .A(fifo_array[426]), .B(n5818), .Y(n625) );
  INVX1 U1429 ( .A(n625), .Y(n3293) );
  AND2X1 U1431 ( .A(fifo_array[405]), .B(n5821), .Y(n603) );
  INVX1 U1433 ( .A(n603), .Y(n3294) );
  AND2X1 U1435 ( .A(fifo_array[396]), .B(n5820), .Y(n594) );
  INVX1 U1437 ( .A(n594), .Y(n3295) );
  AND2X1 U1439 ( .A(fifo_array[383]), .B(n5820), .Y(n581) );
  INVX1 U1441 ( .A(n581), .Y(n3296) );
  AND2X1 U1443 ( .A(fifo_array[353]), .B(n5823), .Y(n549) );
  INVX1 U1445 ( .A(n549), .Y(n3297) );
  AND2X1 U1447 ( .A(fifo_array[340]), .B(n5822), .Y(n536) );
  INVX1 U1449 ( .A(n536), .Y(n3298) );
  AND2X1 U1451 ( .A(fifo_array[324]), .B(n5825), .Y(n518) );
  INVX1 U1453 ( .A(n518), .Y(n3299) );
  AND2X1 U1455 ( .A(fifo_array[318]), .B(n5824), .Y(n512) );
  INVX1 U1457 ( .A(n512), .Y(n3300) );
  AND2X1 U1459 ( .A(fifo_array[306]), .B(n5824), .Y(n500) );
  INVX1 U1461 ( .A(n500), .Y(n3301) );
  AND2X1 U1463 ( .A(fifo_array[291]), .B(n5827), .Y(n483) );
  INVX1 U1465 ( .A(n483), .Y(n3302) );
  AND2X1 U1467 ( .A(fifo_array[275]), .B(n5826), .Y(n467) );
  INVX1 U1469 ( .A(n467), .Y(n3303) );
  AND2X1 U1471 ( .A(fifo_array[263]), .B(n5827), .Y(n455) );
  INVX1 U1473 ( .A(n455), .Y(n3304) );
  AND2X1 U1475 ( .A(fifo_array[246]), .B(n5829), .Y(n436) );
  INVX1 U1477 ( .A(n436), .Y(n3305) );
  AND2X1 U1478 ( .A(fifo_array[232]), .B(n5828), .Y(n422) );
  INVX1 U1481 ( .A(n422), .Y(n3306) );
  AND2X1 U1483 ( .A(fifo_array[220]), .B(n5829), .Y(n410) );
  INVX1 U1485 ( .A(n410), .Y(n3307) );
  AND2X1 U1487 ( .A(fifo_array[184]), .B(n5831), .Y(n372) );
  INVX1 U1489 ( .A(n372), .Y(n3308) );
  AND2X1 U1491 ( .A(fifo_array[177]), .B(n5831), .Y(n365) );
  INVX1 U1493 ( .A(n365), .Y(n3309) );
  AND2X1 U1495 ( .A(fifo_array[166]), .B(n5833), .Y(n352) );
  INVX1 U1497 ( .A(n352), .Y(n3310) );
  AND2X1 U1499 ( .A(fifo_array[160]), .B(n5833), .Y(n346) );
  INVX1 U1501 ( .A(n346), .Y(n3311) );
  AND2X1 U1503 ( .A(fifo_array[117]), .B(n5835), .Y(n301) );
  INVX1 U1505 ( .A(n301), .Y(n3312) );
  AND2X1 U1507 ( .A(fifo_array[80]), .B(n5837), .Y(n262) );
  INVX1 U1509 ( .A(n262), .Y(n3313) );
  AND2X1 U1511 ( .A(fifo_array[74]), .B(n5837), .Y(n256) );
  INVX1 U1513 ( .A(n256), .Y(n3314) );
  AND2X1 U1515 ( .A(fifo_array[37]), .B(n5839), .Y(n216) );
  INVX1 U1517 ( .A(n216), .Y(n3315) );
  AND2X1 U1519 ( .A(fifo_array[31]), .B(n5839), .Y(n210) );
  INVX1 U1521 ( .A(n210), .Y(n3316) );
  AND2X1 U1523 ( .A(fifo_array[1335]), .B(n5776), .Y(n1557) );
  INVX1 U1525 ( .A(n1557), .Y(n3317) );
  AND2X1 U1527 ( .A(fifo_array[1300]), .B(n5779), .Y(n1521) );
  INVX1 U1529 ( .A(n1521), .Y(n3318) );
  AND2X1 U1531 ( .A(fifo_array[1294]), .B(n5778), .Y(n1515) );
  INVX1 U1533 ( .A(n1515), .Y(n3319) );
  AND2X1 U1535 ( .A(fifo_array[1234]), .B(n5781), .Y(n1454) );
  INVX1 U1537 ( .A(n1454), .Y(n3320) );
  AND2X1 U1539 ( .A(fifo_array[1227]), .B(n5780), .Y(n1447) );
  INVX1 U1541 ( .A(n1447), .Y(n3321) );
  AND2X1 U1543 ( .A(fifo_array[1212]), .B(n5783), .Y(n1431) );
  INVX1 U1545 ( .A(n1431), .Y(n3322) );
  AND2X1 U1547 ( .A(fifo_array[1198]), .B(n5782), .Y(n1417) );
  INVX1 U1549 ( .A(n1417), .Y(n3323) );
  AND2X1 U1551 ( .A(fifo_array[1186]), .B(n5782), .Y(n1405) );
  INVX1 U1553 ( .A(n1405), .Y(n3324) );
  AND2X1 U1555 ( .A(fifo_array[1173]), .B(n5785), .Y(n1391) );
  INVX1 U1557 ( .A(n1391), .Y(n3325) );
  AND2X1 U1559 ( .A(fifo_array[1157]), .B(n5784), .Y(n1375) );
  INVX1 U1561 ( .A(n1375), .Y(n3326) );
  AND2X1 U1563 ( .A(fifo_array[1145]), .B(n5784), .Y(n1363) );
  INVX1 U1564 ( .A(n1363), .Y(n3327) );
  AND2X1 U1566 ( .A(fifo_array[1122]), .B(n5786), .Y(n1339) );
  INVX1 U1568 ( .A(n1339), .Y(n3328) );
  AND2X1 U1570 ( .A(fifo_array[1116]), .B(n5786), .Y(n1333) );
  INVX1 U1572 ( .A(n1333), .Y(n3329) );
  AND2X1 U1574 ( .A(fifo_array[1104]), .B(n5787), .Y(n1321) );
  INVX1 U1576 ( .A(n1321), .Y(n3330) );
  AND2X1 U1578 ( .A(fifo_array[1079]), .B(n5788), .Y(n1295) );
  INVX1 U1580 ( .A(n1295), .Y(n3331) );
  AND2X1 U1582 ( .A(fifo_array[1070]), .B(n5789), .Y(n1286) );
  INVX1 U1584 ( .A(n1286), .Y(n3332) );
  AND2X1 U1586 ( .A(fifo_array[1057]), .B(n5789), .Y(n1273) );
  INVX1 U1588 ( .A(n1273), .Y(n3333) );
  AND2X1 U1590 ( .A(fifo_array[1029]), .B(n5791), .Y(n1243) );
  INVX1 U1592 ( .A(n1243), .Y(n3334) );
  AND2X1 U1594 ( .A(fifo_array[1016]), .B(n5790), .Y(n1230) );
  INVX1 U1596 ( .A(n1230), .Y(n3335) );
  AND2X1 U1598 ( .A(fifo_array[1008]), .B(n5791), .Y(n1222) );
  INVX1 U1600 ( .A(n1222), .Y(n3336) );
  AND2X1 U1602 ( .A(fifo_array[991]), .B(n5792), .Y(n1204) );
  INVX1 U1604 ( .A(n1204), .Y(n3337) );
  AND2X1 U1606 ( .A(fifo_array[979]), .B(n5793), .Y(n1192) );
  INVX1 U1608 ( .A(n1192), .Y(n3338) );
  AND2X1 U1610 ( .A(fifo_array[967]), .B(n5793), .Y(n1180) );
  INVX1 U1612 ( .A(n1180), .Y(n3339) );
  AND2X1 U1614 ( .A(fifo_array[950]), .B(n5794), .Y(n1162) );
  INVX1 U1616 ( .A(n1162), .Y(n3340) );
  AND2X1 U1618 ( .A(fifo_array[938]), .B(n5795), .Y(n1150) );
  INVX1 U1620 ( .A(n1150), .Y(n3341) );
  AND2X1 U1622 ( .A(fifo_array[926]), .B(n5795), .Y(n1138) );
  INVX1 U1624 ( .A(n1138), .Y(n3342) );
  AND2X1 U1626 ( .A(fifo_array[897]), .B(n5797), .Y(n1108) );
  INVX1 U1628 ( .A(n1108), .Y(n3343) );
  AND2X1 U1630 ( .A(fifo_array[885]), .B(n5797), .Y(n1096) );
  INVX1 U1632 ( .A(n1096), .Y(n3344) );
  AND2X1 U1634 ( .A(fifo_array[877]), .B(n5798), .Y(n1087) );
  INVX1 U1636 ( .A(n1087), .Y(n3345) );
  AND2X1 U1638 ( .A(fifo_array[871]), .B(n5799), .Y(n1081) );
  INVX1 U1640 ( .A(n1081), .Y(n3346) );
  AND2X1 U1642 ( .A(fifo_array[836]), .B(n5800), .Y(n1045) );
  INVX1 U1644 ( .A(n1045), .Y(n3347) );
  AND2X1 U1646 ( .A(fifo_array[830]), .B(n5801), .Y(n1039) );
  INVX1 U1648 ( .A(n1039), .Y(n3348) );
  AND2X1 U1649 ( .A(fifo_array[789]), .B(n5803), .Y(n997) );
  INVX1 U1651 ( .A(n997), .Y(n3349) );
  AND2X1 U1653 ( .A(fifo_array[754]), .B(n5804), .Y(n961) );
  INVX1 U1655 ( .A(n961), .Y(n3350) );
  AND2X1 U1657 ( .A(fifo_array[748]), .B(n5805), .Y(n955) );
  INVX1 U1659 ( .A(n955), .Y(n3351) );
  AND2X1 U1661 ( .A(fifo_array[688]), .B(n5806), .Y(n893) );
  INVX1 U1663 ( .A(n893), .Y(n3352) );
  AND2X1 U1665 ( .A(fifo_array[681]), .B(n5807), .Y(n886) );
  INVX1 U1667 ( .A(n886), .Y(n3353) );
  AND2X1 U1669 ( .A(fifo_array[666]), .B(n5808), .Y(n870) );
  INVX1 U1671 ( .A(n870), .Y(n3354) );
  AND2X1 U1673 ( .A(fifo_array[652]), .B(n5808), .Y(n856) );
  INVX1 U1675 ( .A(n856), .Y(n3355) );
  AND2X1 U1677 ( .A(fifo_array[640]), .B(n5809), .Y(n844) );
  INVX1 U1679 ( .A(n844), .Y(n3356) );
  AND2X1 U1681 ( .A(fifo_array[627]), .B(n5810), .Y(n830) );
  INVX1 U1683 ( .A(n830), .Y(n3357) );
  AND2X1 U1685 ( .A(fifo_array[611]), .B(n5810), .Y(n814) );
  INVX1 U1687 ( .A(n814), .Y(n3358) );
  AND2X1 U1689 ( .A(fifo_array[599]), .B(n5811), .Y(n802) );
  INVX1 U1691 ( .A(n802), .Y(n3359) );
  AND2X1 U1693 ( .A(fifo_array[576]), .B(n5813), .Y(n778) );
  INVX1 U1695 ( .A(n778), .Y(n3360) );
  AND2X1 U1697 ( .A(fifo_array[570]), .B(n5812), .Y(n772) );
  INVX1 U1699 ( .A(n772), .Y(n3361) );
  AND2X1 U1701 ( .A(fifo_array[558]), .B(n5812), .Y(n760) );
  INVX1 U1703 ( .A(n760), .Y(n3362) );
  AND2X1 U1705 ( .A(fifo_array[533]), .B(n5815), .Y(n734) );
  INVX1 U1707 ( .A(n734), .Y(n3363) );
  AND2X1 U1709 ( .A(fifo_array[524]), .B(n5814), .Y(n725) );
  INVX1 U1711 ( .A(n725), .Y(n3364) );
  AND2X1 U1713 ( .A(fifo_array[511]), .B(n5814), .Y(n712) );
  INVX1 U1715 ( .A(n712), .Y(n3365) );
  AND2X1 U1717 ( .A(fifo_array[483]), .B(n5816), .Y(n683) );
  INVX1 U1719 ( .A(n683), .Y(n3366) );
  AND2X1 U1721 ( .A(fifo_array[470]), .B(n5817), .Y(n670) );
  INVX1 U1723 ( .A(n670), .Y(n3367) );
  AND2X1 U1725 ( .A(fifo_array[462]), .B(n5817), .Y(n662) );
  INVX1 U1727 ( .A(n662), .Y(n3368) );
  AND2X1 U1729 ( .A(fifo_array[445]), .B(n5818), .Y(n644) );
  INVX1 U1731 ( .A(n644), .Y(n3369) );
  AND2X1 U1733 ( .A(fifo_array[433]), .B(n5819), .Y(n632) );
  INVX1 U1734 ( .A(n632), .Y(n3370) );
  AND2X1 U1736 ( .A(fifo_array[421]), .B(n5819), .Y(n620) );
  INVX1 U1738 ( .A(n620), .Y(n3371) );
  AND2X1 U1740 ( .A(fifo_array[404]), .B(n5820), .Y(n602) );
  INVX1 U1742 ( .A(n602), .Y(n3372) );
  AND2X1 U1744 ( .A(fifo_array[392]), .B(n5821), .Y(n590) );
  INVX1 U1746 ( .A(n590), .Y(n3373) );
  AND2X1 U1748 ( .A(fifo_array[380]), .B(n5821), .Y(n578) );
  INVX1 U1750 ( .A(n578), .Y(n3374) );
  AND2X1 U1752 ( .A(fifo_array[351]), .B(n5823), .Y(n547) );
  INVX1 U1754 ( .A(n547), .Y(n3375) );
  AND2X1 U1756 ( .A(fifo_array[339]), .B(n5823), .Y(n535) );
  INVX1 U1758 ( .A(n535), .Y(n3376) );
  AND2X1 U1760 ( .A(fifo_array[331]), .B(n5824), .Y(n525) );
  INVX1 U1762 ( .A(n525), .Y(n3377) );
  AND2X1 U1764 ( .A(fifo_array[325]), .B(n5825), .Y(n519) );
  INVX1 U1766 ( .A(n519), .Y(n3378) );
  AND2X1 U1768 ( .A(fifo_array[290]), .B(n5826), .Y(n482) );
  INVX1 U1770 ( .A(n482), .Y(n3379) );
  AND2X1 U1772 ( .A(fifo_array[284]), .B(n5827), .Y(n476) );
  INVX1 U1774 ( .A(n476), .Y(n3380) );
  AND2X1 U1776 ( .A(fifo_array[243]), .B(n5829), .Y(n433) );
  INVX1 U1778 ( .A(n433), .Y(n3381) );
  AND2X1 U1780 ( .A(fifo_array[208]), .B(n5830), .Y(n396) );
  INVX1 U1782 ( .A(n396), .Y(n3382) );
  AND2X1 U1784 ( .A(fifo_array[202]), .B(n5831), .Y(n390) );
  INVX1 U1786 ( .A(n390), .Y(n3383) );
  AND2X1 U1788 ( .A(fifo_array[142]), .B(n5832), .Y(n328) );
  INVX1 U1790 ( .A(n328), .Y(n3384) );
  AND2X1 U1792 ( .A(fifo_array[135]), .B(n5833), .Y(n321) );
  INVX1 U1794 ( .A(n321), .Y(n3385) );
  AND2X1 U1796 ( .A(fifo_array[120]), .B(n5834), .Y(n304) );
  INVX1 U1798 ( .A(n304), .Y(n3386) );
  AND2X1 U1800 ( .A(fifo_array[106]), .B(n5834), .Y(n290) );
  INVX1 U1802 ( .A(n290), .Y(n3387) );
  AND2X1 U1804 ( .A(fifo_array[94]), .B(n5835), .Y(n278) );
  INVX1 U1806 ( .A(n278), .Y(n3388) );
  AND2X1 U1808 ( .A(fifo_array[81]), .B(n5836), .Y(n263) );
  INVX1 U1810 ( .A(n263), .Y(n3389) );
  AND2X1 U1812 ( .A(fifo_array[65]), .B(n5836), .Y(n247) );
  INVX1 U1814 ( .A(n247), .Y(n3390) );
  AND2X1 U1816 ( .A(fifo_array[53]), .B(n5837), .Y(n235) );
  INVX1 U1818 ( .A(n235), .Y(n3391) );
  AND2X1 U1819 ( .A(fifo_array[30]), .B(n5838), .Y(n209) );
  INVX1 U1821 ( .A(n209), .Y(n3392) );
  AND2X1 U1823 ( .A(fifo_array[24]), .B(n5839), .Y(n203) );
  INVX1 U1825 ( .A(n203), .Y(n3393) );
  AND2X1 U1827 ( .A(fifo_array[12]), .B(n5839), .Y(n191) );
  INVX1 U1829 ( .A(n191), .Y(n3394) );
  AND2X1 U1831 ( .A(fifo_array[1342]), .B(n5777), .Y(n1564) );
  INVX1 U1833 ( .A(n1564), .Y(n3395) );
  AND2X1 U1835 ( .A(fifo_array[1336]), .B(n5776), .Y(n1558) );
  INVX1 U1837 ( .A(n1558), .Y(n3396) );
  AND2X1 U1839 ( .A(fifo_array[1293]), .B(n5778), .Y(n1514) );
  INVX1 U1841 ( .A(n1514), .Y(n3397) );
  AND2X1 U1843 ( .A(fifo_array[1254]), .B(n5781), .Y(n1474) );
  INVX1 U1845 ( .A(n1474), .Y(n3398) );
  AND2X1 U1847 ( .A(fifo_array[1240]), .B(n5780), .Y(n1460) );
  INVX1 U1849 ( .A(n1460), .Y(n3399) );
  AND2X1 U1851 ( .A(fifo_array[1228]), .B(n5780), .Y(n1448) );
  INVX1 U1853 ( .A(n1448), .Y(n3400) );
  AND2X1 U1855 ( .A(fifo_array[1192]), .B(n5783), .Y(n1411) );
  INVX1 U1857 ( .A(n1411), .Y(n3401) );
  AND2X1 U1859 ( .A(fifo_array[1185]), .B(n5782), .Y(n1404) );
  INVX1 U1861 ( .A(n1404), .Y(n3402) );
  AND2X1 U1863 ( .A(fifo_array[1164]), .B(n5784), .Y(n1382) );
  INVX1 U1865 ( .A(n1382), .Y(n3403) );
  AND2X1 U1867 ( .A(fifo_array[1158]), .B(n5785), .Y(n1376) );
  INVX1 U1869 ( .A(n1376), .Y(n3404) );
  AND2X1 U1871 ( .A(fifo_array[1146]), .B(n5785), .Y(n1364) );
  INVX1 U1873 ( .A(n1364), .Y(n3405) );
  AND2X1 U1875 ( .A(fifo_array[1131]), .B(n5787), .Y(n1348) );
  INVX1 U1877 ( .A(n1348), .Y(n3406) );
  AND2X1 U1879 ( .A(fifo_array[1115]), .B(n5787), .Y(n1332) );
  INVX1 U1881 ( .A(n1332), .Y(n3407) );
  AND2X1 U1883 ( .A(fifo_array[1103]), .B(n5786), .Y(n1320) );
  INVX1 U1885 ( .A(n1320), .Y(n3408) );
  AND2X1 U1887 ( .A(fifo_array[1078]), .B(n5789), .Y(n1294) );
  INVX1 U1889 ( .A(n1294), .Y(n3409) );
  AND2X1 U1891 ( .A(fifo_array[1069]), .B(n5789), .Y(n1285) );
  INVX1 U1893 ( .A(n1285), .Y(n3410) );
  AND2X1 U1895 ( .A(fifo_array[1056]), .B(n5789), .Y(n1272) );
  INVX1 U1897 ( .A(n1272), .Y(n3411) );
  AND2X1 U1899 ( .A(fifo_array[1033]), .B(n5791), .Y(n1247) );
  INVX1 U1901 ( .A(n1247), .Y(n3412) );
  AND2X1 U1903 ( .A(fifo_array[1021]), .B(n5791), .Y(n1235) );
  INVX1 U1904 ( .A(n1235), .Y(n3413) );
  AND2X1 U1906 ( .A(fifo_array[1009]), .B(n5791), .Y(n1223) );
  INVX1 U1908 ( .A(n1223), .Y(n3414) );
  AND2X1 U1910 ( .A(fifo_array[987]), .B(n5792), .Y(n1200) );
  INVX1 U1912 ( .A(n1200), .Y(n3415) );
  AND2X1 U1914 ( .A(fifo_array[974]), .B(n5793), .Y(n1187) );
  INVX1 U1916 ( .A(n1187), .Y(n3416) );
  AND2X1 U1918 ( .A(fifo_array[966]), .B(n5793), .Y(n1179) );
  INVX1 U1920 ( .A(n1179), .Y(n3417) );
  AND2X1 U1922 ( .A(fifo_array[939]), .B(n5795), .Y(n1151) );
  INVX1 U1924 ( .A(n1151), .Y(n3418) );
  AND2X1 U1926 ( .A(fifo_array[927]), .B(n5794), .Y(n1139) );
  INVX1 U1928 ( .A(n1139), .Y(n3419) );
  AND2X1 U1930 ( .A(fifo_array[908]), .B(n5796), .Y(n1119) );
  INVX1 U1932 ( .A(n1119), .Y(n3420) );
  AND2X1 U1934 ( .A(fifo_array[896]), .B(n5797), .Y(n1107) );
  INVX1 U1936 ( .A(n1107), .Y(n3421) );
  AND2X1 U1938 ( .A(fifo_array[884]), .B(n5796), .Y(n1095) );
  INVX1 U1940 ( .A(n1095), .Y(n3422) );
  AND2X1 U1942 ( .A(fifo_array[878]), .B(n5799), .Y(n1088) );
  INVX1 U1944 ( .A(n1088), .Y(n3423) );
  AND2X1 U1946 ( .A(fifo_array[872]), .B(n5799), .Y(n1082) );
  INVX1 U1948 ( .A(n1082), .Y(n3424) );
  AND2X1 U1950 ( .A(fifo_array[835]), .B(n5801), .Y(n1044) );
  INVX1 U1952 ( .A(n1044), .Y(n3425) );
  AND2X1 U1954 ( .A(fifo_array[829]), .B(n5801), .Y(n1038) );
  INVX1 U1956 ( .A(n1038), .Y(n3426) );
  AND2X1 U1958 ( .A(fifo_array[796]), .B(n5802), .Y(n1004) );
  INVX1 U1960 ( .A(n1004), .Y(n3427) );
  AND2X1 U1962 ( .A(fifo_array[790]), .B(n5803), .Y(n998) );
  INVX1 U1964 ( .A(n998), .Y(n3428) );
  AND2X1 U1966 ( .A(fifo_array[747]), .B(n5805), .Y(n954) );
  INVX1 U1968 ( .A(n954), .Y(n3429) );
  AND2X1 U1970 ( .A(fifo_array[708]), .B(n5807), .Y(n913) );
  INVX1 U1972 ( .A(n913), .Y(n3430) );
  AND2X1 U1974 ( .A(fifo_array[694]), .B(n5806), .Y(n899) );
  INVX1 U1976 ( .A(n899), .Y(n3431) );
  AND2X1 U1978 ( .A(fifo_array[682]), .B(n5807), .Y(n887) );
  INVX1 U1980 ( .A(n887), .Y(n3432) );
  AND2X1 U1982 ( .A(fifo_array[646]), .B(n5809), .Y(n850) );
  INVX1 U1984 ( .A(n850), .Y(n3433) );
  AND2X1 U1986 ( .A(fifo_array[639]), .B(n5809), .Y(n843) );
  INVX1 U1988 ( .A(n843), .Y(n3434) );
  AND2X1 U1989 ( .A(fifo_array[618]), .B(n5811), .Y(n821) );
  INVX1 U1991 ( .A(n821), .Y(n3435) );
  AND2X1 U1993 ( .A(fifo_array[612]), .B(n5810), .Y(n815) );
  INVX1 U1995 ( .A(n815), .Y(n3436) );
  AND2X1 U1997 ( .A(fifo_array[600]), .B(n5810), .Y(n803) );
  INVX1 U1999 ( .A(n803), .Y(n3437) );
  AND2X1 U2001 ( .A(fifo_array[585]), .B(n5812), .Y(n787) );
  INVX1 U2003 ( .A(n787), .Y(n3438) );
  AND2X1 U2005 ( .A(fifo_array[569]), .B(n5812), .Y(n771) );
  INVX1 U2007 ( .A(n771), .Y(n3439) );
  AND2X1 U2009 ( .A(fifo_array[557]), .B(n5813), .Y(n759) );
  INVX1 U2011 ( .A(n759), .Y(n3440) );
  AND2X1 U2013 ( .A(fifo_array[532]), .B(n5815), .Y(n733) );
  INVX1 U2015 ( .A(n733), .Y(n3441) );
  AND2X1 U2017 ( .A(fifo_array[523]), .B(n5814), .Y(n724) );
  INVX1 U2019 ( .A(n724), .Y(n3442) );
  AND2X1 U2021 ( .A(fifo_array[510]), .B(n5814), .Y(n711) );
  INVX1 U2023 ( .A(n711), .Y(n3443) );
  AND2X1 U2025 ( .A(fifo_array[487]), .B(n5816), .Y(n687) );
  INVX1 U2027 ( .A(n687), .Y(n3444) );
  AND2X1 U2029 ( .A(fifo_array[475]), .B(n5817), .Y(n675) );
  INVX1 U2031 ( .A(n675), .Y(n3445) );
  AND2X1 U2033 ( .A(fifo_array[463]), .B(n5817), .Y(n663) );
  INVX1 U2035 ( .A(n663), .Y(n3446) );
  AND2X1 U2037 ( .A(fifo_array[441]), .B(n5818), .Y(n640) );
  INVX1 U2039 ( .A(n640), .Y(n3447) );
  AND2X1 U2041 ( .A(fifo_array[428]), .B(n5819), .Y(n627) );
  INVX1 U2043 ( .A(n627), .Y(n3448) );
  AND2X1 U2045 ( .A(fifo_array[420]), .B(n5819), .Y(n619) );
  INVX1 U2047 ( .A(n619), .Y(n3449) );
  AND2X1 U2049 ( .A(fifo_array[393]), .B(n5821), .Y(n591) );
  INVX1 U2051 ( .A(n591), .Y(n3450) );
  AND2X1 U2053 ( .A(fifo_array[381]), .B(n5820), .Y(n579) );
  INVX1 U2055 ( .A(n579), .Y(n3451) );
  AND2X1 U2057 ( .A(fifo_array[362]), .B(n5822), .Y(n558) );
  INVX1 U2059 ( .A(n558), .Y(n3452) );
  AND2X1 U2061 ( .A(fifo_array[350]), .B(n5823), .Y(n546) );
  INVX1 U2063 ( .A(n546), .Y(n3453) );
  AND2X1 U2065 ( .A(fifo_array[338]), .B(n5822), .Y(n534) );
  INVX1 U2067 ( .A(n534), .Y(n3454) );
  AND2X1 U2069 ( .A(fifo_array[332]), .B(n5825), .Y(n526) );
  INVX1 U2071 ( .A(n526), .Y(n3455) );
  AND2X1 U2073 ( .A(fifo_array[326]), .B(n5825), .Y(n520) );
  INVX1 U2074 ( .A(n520), .Y(n3456) );
  AND2X1 U2076 ( .A(fifo_array[289]), .B(n5827), .Y(n481) );
  INVX1 U2078 ( .A(n481), .Y(n3457) );
  AND2X1 U2080 ( .A(fifo_array[283]), .B(n5827), .Y(n475) );
  INVX1 U2082 ( .A(n475), .Y(n3458) );
  AND2X1 U2084 ( .A(fifo_array[250]), .B(n5828), .Y(n440) );
  INVX1 U2086 ( .A(n440), .Y(n3459) );
  AND2X1 U2088 ( .A(fifo_array[244]), .B(n5829), .Y(n434) );
  INVX1 U2090 ( .A(n434), .Y(n3460) );
  AND2X1 U2092 ( .A(fifo_array[201]), .B(n5831), .Y(n389) );
  INVX1 U2094 ( .A(n389), .Y(n3461) );
  AND2X1 U2096 ( .A(fifo_array[162]), .B(n5833), .Y(n348) );
  INVX1 U2098 ( .A(n348), .Y(n3462) );
  AND2X1 U2100 ( .A(fifo_array[148]), .B(n5832), .Y(n334) );
  INVX1 U2102 ( .A(n334), .Y(n3463) );
  AND2X1 U2104 ( .A(fifo_array[136]), .B(n5833), .Y(n322) );
  INVX1 U2106 ( .A(n322), .Y(n3464) );
  AND2X1 U2108 ( .A(fifo_array[100]), .B(n5835), .Y(n284) );
  INVX1 U2110 ( .A(n284), .Y(n3465) );
  AND2X1 U2112 ( .A(fifo_array[93]), .B(n5835), .Y(n277) );
  INVX1 U2114 ( .A(n277), .Y(n3466) );
  AND2X1 U2116 ( .A(fifo_array[72]), .B(n5837), .Y(n254) );
  INVX1 U2118 ( .A(n254), .Y(n3467) );
  AND2X1 U2120 ( .A(fifo_array[66]), .B(n5836), .Y(n248) );
  INVX1 U2122 ( .A(n248), .Y(n3468) );
  AND2X1 U2124 ( .A(fifo_array[54]), .B(n5836), .Y(n236) );
  INVX1 U2126 ( .A(n236), .Y(n3469) );
  AND2X1 U2128 ( .A(fifo_array[39]), .B(n5839), .Y(n218) );
  INVX1 U2130 ( .A(n218), .Y(n3470) );
  AND2X1 U2132 ( .A(fifo_array[23]), .B(n5839), .Y(n202) );
  INVX1 U2134 ( .A(n202), .Y(n3471) );
  AND2X1 U2136 ( .A(fifo_array[11]), .B(n5839), .Y(n190) );
  INVX1 U2138 ( .A(n190), .Y(n3472) );
  AND2X1 U2140 ( .A(fifo_array[1339]), .B(n5777), .Y(n1561) );
  INVX1 U2142 ( .A(n1561), .Y(n3473) );
  AND2X1 U2144 ( .A(fifo_array[1333]), .B(n5776), .Y(n1555) );
  INVX1 U2146 ( .A(n1555), .Y(n3474) );
  AND2X1 U2148 ( .A(fifo_array[1298]), .B(n5779), .Y(n1519) );
  INVX1 U2150 ( .A(n1519), .Y(n3475) );
  AND2X1 U2152 ( .A(fifo_array[1292]), .B(n5778), .Y(n1513) );
  INVX1 U2154 ( .A(n1513), .Y(n3476) );
  AND2X1 U2156 ( .A(fifo_array[1257]), .B(n5781), .Y(n1477) );
  INVX1 U2158 ( .A(n1477), .Y(n3477) );
  AND2X1 U2159 ( .A(fifo_array[1241]), .B(n5781), .Y(n1461) );
  INVX1 U2162 ( .A(n1461), .Y(n3478) );
  AND2X1 U2164 ( .A(fifo_array[1229]), .B(n5780), .Y(n1449) );
  INVX1 U2166 ( .A(n1449), .Y(n3479) );
  AND2X1 U2168 ( .A(fifo_array[1206]), .B(n5782), .Y(n1425) );
  INVX1 U2170 ( .A(n1425), .Y(n3480) );
  AND2X1 U2172 ( .A(fifo_array[1200]), .B(n5783), .Y(n1419) );
  INVX1 U2174 ( .A(n1419), .Y(n3481) );
  AND2X1 U2176 ( .A(fifo_array[1188]), .B(n5783), .Y(n1407) );
  INVX1 U2178 ( .A(n1407), .Y(n3482) );
  AND2X1 U2180 ( .A(fifo_array[1150]), .B(n5785), .Y(n1368) );
  INVX1 U2182 ( .A(n1368), .Y(n3483) );
  AND2X1 U2184 ( .A(fifo_array[1143]), .B(n5784), .Y(n1361) );
  INVX1 U2186 ( .A(n1361), .Y(n3484) );
  AND2X1 U2188 ( .A(fifo_array[1128]), .B(n5787), .Y(n1345) );
  INVX1 U2190 ( .A(n1345), .Y(n3485) );
  AND2X1 U2192 ( .A(fifo_array[1114]), .B(n5786), .Y(n1331) );
  INVX1 U2194 ( .A(n1331), .Y(n3486) );
  AND2X1 U2196 ( .A(fifo_array[1102]), .B(n5786), .Y(n1319) );
  INVX1 U2198 ( .A(n1319), .Y(n3487) );
  AND2X1 U2200 ( .A(fifo_array[1077]), .B(n5788), .Y(n1293) );
  INVX1 U2202 ( .A(n1293), .Y(n3488) );
  AND2X1 U2204 ( .A(fifo_array[1068]), .B(n5788), .Y(n1284) );
  INVX1 U2206 ( .A(n1284), .Y(n3489) );
  AND2X1 U2208 ( .A(fifo_array[1055]), .B(n5789), .Y(n1271) );
  INVX1 U2210 ( .A(n1271), .Y(n3490) );
  AND2X1 U2212 ( .A(fifo_array[1034]), .B(n5790), .Y(n1248) );
  INVX1 U2214 ( .A(n1248), .Y(n3491) );
  AND2X1 U2216 ( .A(fifo_array[1022]), .B(n5791), .Y(n1236) );
  INVX1 U2218 ( .A(n1236), .Y(n3492) );
  AND2X1 U2220 ( .A(fifo_array[1010]), .B(n5791), .Y(n1224) );
  INVX1 U2222 ( .A(n1224), .Y(n3493) );
  AND2X1 U2224 ( .A(fifo_array[981]), .B(n5793), .Y(n1194) );
  INVX1 U2226 ( .A(n1194), .Y(n3494) );
  AND2X1 U2228 ( .A(fifo_array[969]), .B(n5793), .Y(n1182) );
  INVX1 U2230 ( .A(n1182), .Y(n3495) );
  AND2X1 U2232 ( .A(fifo_array[945]), .B(n5794), .Y(n1157) );
  INVX1 U2234 ( .A(n1157), .Y(n3496) );
  AND2X1 U2236 ( .A(fifo_array[932]), .B(n5795), .Y(n1144) );
  INVX1 U2238 ( .A(n1144), .Y(n3497) );
  AND2X1 U2240 ( .A(fifo_array[924]), .B(n5795), .Y(n1136) );
  INVX1 U2242 ( .A(n1136), .Y(n3498) );
  AND2X1 U2244 ( .A(fifo_array[907]), .B(n5796), .Y(n1118) );
  INVX1 U2245 ( .A(n1118), .Y(n3499) );
  AND2X1 U2248 ( .A(fifo_array[895]), .B(n5797), .Y(n1106) );
  INVX1 U2250 ( .A(n1106), .Y(n3500) );
  AND2X1 U2252 ( .A(fifo_array[883]), .B(n5797), .Y(n1094) );
  INVX1 U2254 ( .A(n1094), .Y(n3501) );
  AND2X1 U2256 ( .A(fifo_array[873]), .B(n5799), .Y(n1083) );
  INVX1 U2258 ( .A(n1083), .Y(n3502) );
  AND2X1 U2260 ( .A(fifo_array[838]), .B(n5800), .Y(n1047) );
  INVX1 U2262 ( .A(n1047), .Y(n3503) );
  AND2X1 U2264 ( .A(fifo_array[832]), .B(n5801), .Y(n1041) );
  INVX1 U2266 ( .A(n1041), .Y(n3504) );
  AND2X1 U2268 ( .A(fifo_array[793]), .B(n5803), .Y(n1001) );
  INVX1 U2270 ( .A(n1001), .Y(n3505) );
  AND2X1 U2272 ( .A(fifo_array[787]), .B(n5803), .Y(n995) );
  INVX1 U2274 ( .A(n995), .Y(n3506) );
  AND2X1 U2276 ( .A(fifo_array[752]), .B(n5805), .Y(n959) );
  INVX1 U2278 ( .A(n959), .Y(n3507) );
  AND2X1 U2280 ( .A(fifo_array[746]), .B(n5805), .Y(n953) );
  INVX1 U2282 ( .A(n953), .Y(n3508) );
  AND2X1 U2284 ( .A(fifo_array[711]), .B(n5806), .Y(n916) );
  INVX1 U2286 ( .A(n916), .Y(n3509) );
  AND2X1 U2288 ( .A(fifo_array[695]), .B(n5806), .Y(n900) );
  INVX1 U2290 ( .A(n900), .Y(n3510) );
  AND2X1 U2292 ( .A(fifo_array[683]), .B(n5807), .Y(n888) );
  INVX1 U2294 ( .A(n888), .Y(n3511) );
  AND2X1 U2296 ( .A(fifo_array[660]), .B(n5809), .Y(n864) );
  INVX1 U2298 ( .A(n864), .Y(n3512) );
  AND2X1 U2300 ( .A(fifo_array[654]), .B(n5808), .Y(n858) );
  INVX1 U2302 ( .A(n858), .Y(n3513) );
  AND2X1 U2304 ( .A(fifo_array[642]), .B(n5808), .Y(n846) );
  INVX1 U2306 ( .A(n846), .Y(n3514) );
  AND2X1 U2308 ( .A(fifo_array[604]), .B(n5811), .Y(n807) );
  INVX1 U2310 ( .A(n807), .Y(n3515) );
  AND2X1 U2312 ( .A(fifo_array[597]), .B(n5811), .Y(n800) );
  INVX1 U2314 ( .A(n800), .Y(n3516) );
  AND2X1 U2316 ( .A(fifo_array[582]), .B(n5813), .Y(n784) );
  INVX1 U2318 ( .A(n784), .Y(n3517) );
  AND2X1 U2320 ( .A(fifo_array[568]), .B(n5812), .Y(n770) );
  INVX1 U2322 ( .A(n770), .Y(n3518) );
  AND2X1 U2324 ( .A(fifo_array[556]), .B(n5813), .Y(n758) );
  INVX1 U2326 ( .A(n758), .Y(n3519) );
  AND2X1 U2328 ( .A(fifo_array[531]), .B(n5815), .Y(n732) );
  INVX1 U2330 ( .A(n732), .Y(n3520) );
  AND2X1 U2331 ( .A(fifo_array[522]), .B(n5814), .Y(n723) );
  INVX1 U2334 ( .A(n723), .Y(n3521) );
  AND2X1 U2336 ( .A(fifo_array[509]), .B(n5815), .Y(n710) );
  INVX1 U2338 ( .A(n710), .Y(n3522) );
  AND2X1 U2340 ( .A(fifo_array[488]), .B(n5816), .Y(n688) );
  INVX1 U2342 ( .A(n688), .Y(n3523) );
  AND2X1 U2344 ( .A(fifo_array[476]), .B(n5817), .Y(n676) );
  INVX1 U2346 ( .A(n676), .Y(n3524) );
  AND2X1 U2348 ( .A(fifo_array[464]), .B(n5817), .Y(n664) );
  INVX1 U2350 ( .A(n664), .Y(n3525) );
  AND2X1 U2352 ( .A(fifo_array[435]), .B(n5819), .Y(n634) );
  INVX1 U2354 ( .A(n634), .Y(n3526) );
  AND2X1 U2356 ( .A(fifo_array[423]), .B(n5819), .Y(n622) );
  INVX1 U2358 ( .A(n622), .Y(n3527) );
  AND2X1 U2360 ( .A(fifo_array[399]), .B(n5820), .Y(n597) );
  INVX1 U2362 ( .A(n597), .Y(n3528) );
  AND2X1 U2364 ( .A(fifo_array[386]), .B(n5821), .Y(n584) );
  INVX1 U2366 ( .A(n584), .Y(n3529) );
  AND2X1 U2368 ( .A(fifo_array[378]), .B(n5821), .Y(n576) );
  INVX1 U2370 ( .A(n576), .Y(n3530) );
  AND2X1 U2372 ( .A(fifo_array[361]), .B(n5822), .Y(n557) );
  INVX1 U2374 ( .A(n557), .Y(n3531) );
  AND2X1 U2376 ( .A(fifo_array[349]), .B(n5823), .Y(n545) );
  INVX1 U2378 ( .A(n545), .Y(n3532) );
  AND2X1 U2380 ( .A(fifo_array[337]), .B(n5823), .Y(n533) );
  INVX1 U2382 ( .A(n533), .Y(n3533) );
  AND2X1 U2384 ( .A(fifo_array[327]), .B(n5825), .Y(n521) );
  INVX1 U2386 ( .A(n521), .Y(n3534) );
  AND2X1 U2388 ( .A(fifo_array[292]), .B(n5826), .Y(n484) );
  INVX1 U2390 ( .A(n484), .Y(n3535) );
  AND2X1 U2392 ( .A(fifo_array[286]), .B(n5827), .Y(n478) );
  INVX1 U2394 ( .A(n478), .Y(n3536) );
  AND2X1 U2396 ( .A(fifo_array[247]), .B(n5829), .Y(n437) );
  INVX1 U2398 ( .A(n437), .Y(n3537) );
  AND2X1 U2400 ( .A(fifo_array[241]), .B(n5829), .Y(n431) );
  INVX1 U2402 ( .A(n431), .Y(n3538) );
  AND2X1 U2404 ( .A(fifo_array[206]), .B(n5831), .Y(n394) );
  INVX1 U2406 ( .A(n394), .Y(n3539) );
  AND2X1 U2408 ( .A(fifo_array[200]), .B(n5831), .Y(n388) );
  INVX1 U2410 ( .A(n388), .Y(n3540) );
  AND2X1 U2412 ( .A(fifo_array[165]), .B(n5832), .Y(n351) );
  INVX1 U2414 ( .A(n351), .Y(n3541) );
  AND2X1 U2416 ( .A(fifo_array[149]), .B(n5832), .Y(n335) );
  INVX1 U2417 ( .A(n335), .Y(n3542) );
  AND2X1 U2420 ( .A(fifo_array[137]), .B(n5833), .Y(n323) );
  INVX1 U2422 ( .A(n323), .Y(n3543) );
  AND2X1 U2424 ( .A(fifo_array[114]), .B(n5835), .Y(n298) );
  INVX1 U2426 ( .A(n298), .Y(n3544) );
  AND2X1 U2428 ( .A(fifo_array[108]), .B(n5834), .Y(n292) );
  INVX1 U2430 ( .A(n292), .Y(n3545) );
  AND2X1 U2432 ( .A(fifo_array[96]), .B(n5834), .Y(n280) );
  INVX1 U2434 ( .A(n280), .Y(n3546) );
  AND2X1 U2436 ( .A(fifo_array[58]), .B(n5837), .Y(n240) );
  INVX1 U2438 ( .A(n240), .Y(n3547) );
  AND2X1 U2440 ( .A(fifo_array[51]), .B(n5837), .Y(n233) );
  INVX1 U2442 ( .A(n233), .Y(n3548) );
  AND2X1 U2444 ( .A(fifo_array[36]), .B(n5839), .Y(n215) );
  INVX1 U2446 ( .A(n215), .Y(n3549) );
  AND2X1 U2448 ( .A(fifo_array[22]), .B(n5839), .Y(n201) );
  INVX1 U2450 ( .A(n201), .Y(n3550) );
  AND2X1 U2452 ( .A(fifo_array[10]), .B(n5838), .Y(n189) );
  INVX1 U2454 ( .A(n189), .Y(n3551) );
  AND2X1 U2456 ( .A(fifo_array[1340]), .B(n5777), .Y(n1562) );
  INVX1 U2458 ( .A(n1562), .Y(n3552) );
  AND2X1 U2460 ( .A(fifo_array[1334]), .B(n5776), .Y(n1556) );
  INVX1 U2462 ( .A(n1556), .Y(n3553) );
  AND2X1 U2464 ( .A(fifo_array[1297]), .B(n5779), .Y(n1518) );
  INVX1 U2466 ( .A(n1518), .Y(n3554) );
  AND2X1 U2468 ( .A(fifo_array[1291]), .B(n5778), .Y(n1512) );
  INVX1 U2470 ( .A(n1512), .Y(n3555) );
  AND2X1 U2472 ( .A(fifo_array[1248]), .B(n5780), .Y(n1468) );
  INVX1 U2474 ( .A(n1468), .Y(n3556) );
  AND2X1 U2476 ( .A(fifo_array[1242]), .B(n5780), .Y(n1462) );
  INVX1 U2478 ( .A(n1462), .Y(n3557) );
  AND2X1 U2480 ( .A(fifo_array[1230]), .B(n5781), .Y(n1450) );
  INVX1 U2482 ( .A(n1450), .Y(n3558) );
  AND2X1 U2484 ( .A(fifo_array[1215]), .B(n5783), .Y(n1434) );
  INVX1 U2486 ( .A(n1434), .Y(n3559) );
  AND2X1 U2488 ( .A(fifo_array[1199]), .B(n5782), .Y(n1418) );
  INVX1 U2490 ( .A(n1418), .Y(n3560) );
  AND2X1 U2492 ( .A(fifo_array[1187]), .B(n5782), .Y(n1406) );
  INVX1 U2494 ( .A(n1406), .Y(n3561) );
  AND2X1 U2496 ( .A(fifo_array[1170]), .B(n5785), .Y(n1388) );
  INVX1 U2498 ( .A(n1388), .Y(n3562) );
  AND2X1 U2500 ( .A(fifo_array[1156]), .B(n5784), .Y(n1374) );
  INVX1 U2502 ( .A(n1374), .Y(n3563) );
  AND2X1 U2503 ( .A(fifo_array[1144]), .B(n5784), .Y(n1362) );
  INVX1 U2506 ( .A(n1362), .Y(n3564) );
  AND2X1 U2508 ( .A(fifo_array[1108]), .B(n5787), .Y(n1325) );
  INVX1 U2510 ( .A(n1325), .Y(n3565) );
  AND2X1 U2512 ( .A(fifo_array[1101]), .B(n5786), .Y(n1318) );
  INVX1 U2514 ( .A(n1318), .Y(n3566) );
  AND2X1 U2516 ( .A(fifo_array[1067]), .B(n5789), .Y(n1283) );
  INVX1 U2518 ( .A(n1283), .Y(n3567) );
  AND2X1 U2520 ( .A(fifo_array[1054]), .B(n5789), .Y(n1270) );
  INVX1 U2522 ( .A(n1270), .Y(n3568) );
  AND2X1 U2524 ( .A(fifo_array[1023]), .B(n5790), .Y(n1237) );
  INVX1 U2526 ( .A(n1237), .Y(n3569) );
  AND2X1 U2528 ( .A(fifo_array[1011]), .B(n5791), .Y(n1225) );
  INVX1 U2530 ( .A(n1225), .Y(n3570) );
  AND2X1 U2532 ( .A(fifo_array[992]), .B(n5792), .Y(n1205) );
  INVX1 U2534 ( .A(n1205), .Y(n3571) );
  AND2X1 U2536 ( .A(fifo_array[980]), .B(n5793), .Y(n1193) );
  INVX1 U2538 ( .A(n1193), .Y(n3572) );
  AND2X1 U2540 ( .A(fifo_array[968]), .B(n5792), .Y(n1181) );
  INVX1 U2542 ( .A(n1181), .Y(n3573) );
  AND2X1 U2544 ( .A(fifo_array[949]), .B(n5794), .Y(n1161) );
  INVX1 U2546 ( .A(n1161), .Y(n3574) );
  AND2X1 U2548 ( .A(fifo_array[937]), .B(n5795), .Y(n1149) );
  INVX1 U2550 ( .A(n1149), .Y(n3575) );
  AND2X1 U2552 ( .A(fifo_array[925]), .B(n5795), .Y(n1137) );
  INVX1 U2554 ( .A(n1137), .Y(n3576) );
  AND2X1 U2556 ( .A(fifo_array[903]), .B(n5796), .Y(n1114) );
  INVX1 U2558 ( .A(n1114), .Y(n3577) );
  AND2X1 U2560 ( .A(fifo_array[890]), .B(n5797), .Y(n1101) );
  INVX1 U2562 ( .A(n1101), .Y(n3578) );
  AND2X1 U2564 ( .A(fifo_array[882]), .B(n5797), .Y(n1093) );
  INVX1 U2566 ( .A(n1093), .Y(n3579) );
  AND2X1 U2568 ( .A(fifo_array[880]), .B(n5798), .Y(n1090) );
  INVX1 U2570 ( .A(n1090), .Y(n3580) );
  AND2X1 U2572 ( .A(fifo_array[874]), .B(n5799), .Y(n1084) );
  INVX1 U2574 ( .A(n1084), .Y(n3581) );
  AND2X1 U2576 ( .A(fifo_array[831]), .B(n5801), .Y(n1040) );
  INVX1 U2578 ( .A(n1040), .Y(n3582) );
  AND2X1 U2580 ( .A(fifo_array[794]), .B(n5802), .Y(n1002) );
  INVX1 U2582 ( .A(n1002), .Y(n3583) );
  AND2X1 U2584 ( .A(fifo_array[788]), .B(n5803), .Y(n996) );
  INVX1 U2586 ( .A(n996), .Y(n3584) );
  AND2X1 U2588 ( .A(fifo_array[751]), .B(n5804), .Y(n958) );
  INVX1 U2589 ( .A(n958), .Y(n3585) );
  AND2X1 U2592 ( .A(fifo_array[745]), .B(n5805), .Y(n952) );
  INVX1 U2594 ( .A(n952), .Y(n3586) );
  AND2X1 U2596 ( .A(fifo_array[702]), .B(n5807), .Y(n907) );
  INVX1 U2598 ( .A(n907), .Y(n3587) );
  AND2X1 U2600 ( .A(fifo_array[696]), .B(n5806), .Y(n901) );
  INVX1 U2602 ( .A(n901), .Y(n3588) );
  AND2X1 U2604 ( .A(fifo_array[684]), .B(n5806), .Y(n889) );
  INVX1 U2606 ( .A(n889), .Y(n3589) );
  AND2X1 U2608 ( .A(fifo_array[669]), .B(n5808), .Y(n873) );
  INVX1 U2610 ( .A(n873), .Y(n3590) );
  AND2X1 U2612 ( .A(fifo_array[653]), .B(n5808), .Y(n857) );
  INVX1 U2614 ( .A(n857), .Y(n3591) );
  AND2X1 U2616 ( .A(fifo_array[641]), .B(n5809), .Y(n845) );
  INVX1 U2618 ( .A(n845), .Y(n3592) );
  AND2X1 U2620 ( .A(fifo_array[624]), .B(n5810), .Y(n827) );
  INVX1 U2622 ( .A(n827), .Y(n3593) );
  AND2X1 U2624 ( .A(fifo_array[610]), .B(n5810), .Y(n813) );
  INVX1 U2626 ( .A(n813), .Y(n3594) );
  AND2X1 U2628 ( .A(fifo_array[598]), .B(n5811), .Y(n801) );
  INVX1 U2630 ( .A(n801), .Y(n3595) );
  AND2X1 U2632 ( .A(fifo_array[562]), .B(n5812), .Y(n764) );
  INVX1 U2634 ( .A(n764), .Y(n3596) );
  AND2X1 U2636 ( .A(fifo_array[555]), .B(n5813), .Y(n757) );
  INVX1 U2638 ( .A(n757), .Y(n3597) );
  AND2X1 U2640 ( .A(fifo_array[521]), .B(n5815), .Y(n722) );
  INVX1 U2642 ( .A(n722), .Y(n3598) );
  AND2X1 U2644 ( .A(fifo_array[508]), .B(n5814), .Y(n709) );
  INVX1 U2646 ( .A(n709), .Y(n3599) );
  AND2X1 U2648 ( .A(fifo_array[477]), .B(n5817), .Y(n677) );
  INVX1 U2650 ( .A(n677), .Y(n3600) );
  AND2X1 U2652 ( .A(fifo_array[465]), .B(n5816), .Y(n665) );
  INVX1 U2654 ( .A(n665), .Y(n3601) );
  AND2X1 U2656 ( .A(fifo_array[446]), .B(n5818), .Y(n645) );
  INVX1 U2658 ( .A(n645), .Y(n3602) );
  AND2X1 U2660 ( .A(fifo_array[434]), .B(n5819), .Y(n633) );
  INVX1 U2662 ( .A(n633), .Y(n3603) );
  AND2X1 U2664 ( .A(fifo_array[422]), .B(n5818), .Y(n621) );
  INVX1 U2666 ( .A(n621), .Y(n3604) );
  AND2X1 U2668 ( .A(fifo_array[403]), .B(n5820), .Y(n601) );
  INVX1 U2670 ( .A(n601), .Y(n3605) );
  AND2X1 U2672 ( .A(fifo_array[391]), .B(n5821), .Y(n589) );
  INVX1 U2674 ( .A(n589), .Y(n3606) );
  AND2X1 U2675 ( .A(fifo_array[379]), .B(n5821), .Y(n577) );
  INVX1 U2678 ( .A(n577), .Y(n3607) );
  AND2X1 U2680 ( .A(fifo_array[357]), .B(n5822), .Y(n553) );
  INVX1 U2682 ( .A(n553), .Y(n3608) );
  AND2X1 U2684 ( .A(fifo_array[344]), .B(n5823), .Y(n540) );
  INVX1 U2686 ( .A(n540), .Y(n3609) );
  AND2X1 U2688 ( .A(fifo_array[336]), .B(n5823), .Y(n532) );
  INVX1 U2690 ( .A(n532), .Y(n3610) );
  AND2X1 U2692 ( .A(fifo_array[334]), .B(n5824), .Y(n528) );
  INVX1 U2694 ( .A(n528), .Y(n3611) );
  AND2X1 U2696 ( .A(fifo_array[328]), .B(n5825), .Y(n522) );
  INVX1 U2698 ( .A(n522), .Y(n3612) );
  AND2X1 U2700 ( .A(fifo_array[285]), .B(n5827), .Y(n477) );
  INVX1 U2702 ( .A(n477), .Y(n3613) );
  AND2X1 U2704 ( .A(fifo_array[248]), .B(n5828), .Y(n438) );
  INVX1 U2706 ( .A(n438), .Y(n3614) );
  AND2X1 U2708 ( .A(fifo_array[242]), .B(n5829), .Y(n432) );
  INVX1 U2710 ( .A(n432), .Y(n3615) );
  AND2X1 U2712 ( .A(fifo_array[205]), .B(n5830), .Y(n393) );
  INVX1 U2714 ( .A(n393), .Y(n3616) );
  AND2X1 U2716 ( .A(fifo_array[199]), .B(n5831), .Y(n387) );
  INVX1 U2718 ( .A(n387), .Y(n3617) );
  AND2X1 U2720 ( .A(fifo_array[156]), .B(n5833), .Y(n342) );
  INVX1 U2722 ( .A(n342), .Y(n3618) );
  AND2X1 U2724 ( .A(fifo_array[150]), .B(n5832), .Y(n336) );
  INVX1 U2726 ( .A(n336), .Y(n3619) );
  AND2X1 U2728 ( .A(fifo_array[138]), .B(n5832), .Y(n324) );
  INVX1 U2730 ( .A(n324), .Y(n3620) );
  AND2X1 U2732 ( .A(fifo_array[123]), .B(n5834), .Y(n307) );
  INVX1 U2734 ( .A(n307), .Y(n3621) );
  AND2X1 U2736 ( .A(fifo_array[107]), .B(n5834), .Y(n291) );
  INVX1 U2738 ( .A(n291), .Y(n3622) );
  AND2X1 U2740 ( .A(fifo_array[95]), .B(n5835), .Y(n279) );
  INVX1 U2742 ( .A(n279), .Y(n3623) );
  AND2X1 U2744 ( .A(fifo_array[78]), .B(n5836), .Y(n260) );
  INVX1 U2746 ( .A(n260), .Y(n3624) );
  AND2X1 U2748 ( .A(fifo_array[64]), .B(n5836), .Y(n246) );
  INVX1 U2750 ( .A(n246), .Y(n3625) );
  AND2X1 U2752 ( .A(fifo_array[52]), .B(n5837), .Y(n234) );
  INVX1 U2754 ( .A(n234), .Y(n3626) );
  AND2X1 U2756 ( .A(fifo_array[16]), .B(n5839), .Y(n195) );
  INVX1 U2758 ( .A(n195), .Y(n3627) );
  AND2X1 U2760 ( .A(fifo_array[9]), .B(n5839), .Y(n188) );
  INVX1 U2761 ( .A(n188), .Y(n3628) );
  AND2X1 U2764 ( .A(n5898), .B(n4231), .Y(n1572) );
  INVX1 U2766 ( .A(n1572), .Y(n3629) );
  AND2X1 U2768 ( .A(fifo_array[1328]), .B(n5777), .Y(n1550) );
  INVX1 U2770 ( .A(n1550), .Y(n3630) );
  AND2X1 U2772 ( .A(fifo_array[1316]), .B(n5776), .Y(n1538) );
  INVX1 U2774 ( .A(n1538), .Y(n3631) );
  AND2X1 U2776 ( .A(fifo_array[1304]), .B(n5777), .Y(n1526) );
  INVX1 U2778 ( .A(n1526), .Y(n3632) );
  AND2X1 U2780 ( .A(fifo_array[1275]), .B(n5778), .Y(n1496) );
  INVX1 U2782 ( .A(n1496), .Y(n3633) );
  AND2X1 U2784 ( .A(fifo_array[1263]), .B(n5779), .Y(n1484) );
  INVX1 U2786 ( .A(n1484), .Y(n3634) );
  AND2X1 U2788 ( .A(fifo_array[1235]), .B(n5780), .Y(n1455) );
  INVX1 U2790 ( .A(n1455), .Y(n3635) );
  AND2X1 U2792 ( .A(fifo_array[1222]), .B(n5781), .Y(n1442) );
  INVX1 U2794 ( .A(n1442), .Y(n3636) );
  AND2X1 U2796 ( .A(fifo_array[1203]), .B(n5782), .Y(n1422) );
  INVX1 U2798 ( .A(n1422), .Y(n3637) );
  AND2X1 U2800 ( .A(fifo_array[1194]), .B(n5783), .Y(n1413) );
  INVX1 U2802 ( .A(n1413), .Y(n3638) );
  AND2X1 U2804 ( .A(fifo_array[1181]), .B(n5783), .Y(n1400) );
  INVX1 U2806 ( .A(n1400), .Y(n3639) );
  AND2X1 U2808 ( .A(fifo_array[1162]), .B(n5784), .Y(n1380) );
  INVX1 U2810 ( .A(n1380), .Y(n3640) );
  AND2X1 U2812 ( .A(fifo_array[1153]), .B(n5785), .Y(n1371) );
  INVX1 U2814 ( .A(n1371), .Y(n3641) );
  AND2X1 U2816 ( .A(fifo_array[1140]), .B(n5785), .Y(n1358) );
  INVX1 U2818 ( .A(n1358), .Y(n3642) );
  AND2X1 U2820 ( .A(fifo_array[1121]), .B(n5786), .Y(n1338) );
  INVX1 U2822 ( .A(n1338), .Y(n3643) );
  AND2X1 U2824 ( .A(fifo_array[1112]), .B(n5787), .Y(n1329) );
  INVX1 U2826 ( .A(n1329), .Y(n3644) );
  AND2X1 U2828 ( .A(fifo_array[1099]), .B(n5787), .Y(n1316) );
  INVX1 U2830 ( .A(n1316), .Y(n3645) );
  AND2X1 U2832 ( .A(fifo_array[1080]), .B(n5788), .Y(n1296) );
  INVX1 U2834 ( .A(n1296), .Y(n3646) );
  AND2X1 U2836 ( .A(fifo_array[1074]), .B(n5788), .Y(n1290) );
  INVX1 U2838 ( .A(n1290), .Y(n3647) );
  AND2X1 U2840 ( .A(fifo_array[1062]), .B(n5789), .Y(n1278) );
  INVX1 U2842 ( .A(n1278), .Y(n3648) );
  AND2X1 U2844 ( .A(fifo_array[1045]), .B(n5791), .Y(n1259) );
  INVX1 U2846 ( .A(n1259), .Y(n3649) );
  AND2X1 U2847 ( .A(fifo_array[1039]), .B(n5790), .Y(n1253) );
  INVX1 U2851 ( .A(n1253), .Y(n3650) );
  AND2X1 U2853 ( .A(fifo_array[1004]), .B(n5793), .Y(n1217) );
  INVX1 U2855 ( .A(n1217), .Y(n3651) );
  AND2X1 U2857 ( .A(fifo_array[998]), .B(n5793), .Y(n1211) );
  INVX1 U2859 ( .A(n1211), .Y(n3652) );
  AND2X1 U2860 ( .A(fifo_array[957]), .B(n5795), .Y(n1169) );
  INVX1 U2861 ( .A(n1169), .Y(n3653) );
  AND2X1 U2873 ( .A(fifo_array[922]), .B(n5797), .Y(n1133) );
  INVX1 U2875 ( .A(n1133), .Y(n3654) );
  AND2X1 U2877 ( .A(fifo_array[916]), .B(n5797), .Y(n1127) );
  INVX1 U2879 ( .A(n1127), .Y(n3655) );
  AND2X1 U2881 ( .A(fifo_array[861]), .B(n5798), .Y(n1071) );
  INVX1 U2882 ( .A(n1071), .Y(n3656) );
  AND2X1 U2925 ( .A(fifo_array[848]), .B(n5799), .Y(n1058) );
  INVX1 U2927 ( .A(n1058), .Y(n3657) );
  AND2X1 U2931 ( .A(fifo_array[840]), .B(n5799), .Y(n1050) );
  INVX1 U2934 ( .A(n1050), .Y(n3658) );
  AND2X1 U2936 ( .A(fifo_array[823]), .B(n5800), .Y(n1032) );
  INVX1 U2941 ( .A(n1032), .Y(n3659) );
  AND2X1 U2942 ( .A(fifo_array[811]), .B(n5801), .Y(n1020) );
  INVX1 U2944 ( .A(n1020), .Y(n3660) );
  AND2X1 U2945 ( .A(fifo_array[799]), .B(n5801), .Y(n1008) );
  INVX1 U2946 ( .A(n1008), .Y(n3661) );
  AND2X1 U2947 ( .A(fifo_array[782]), .B(n5802), .Y(n990) );
  INVX1 U2948 ( .A(n990), .Y(n3662) );
  AND2X1 U2949 ( .A(fifo_array[770]), .B(n5803), .Y(n978) );
  INVX1 U2950 ( .A(n978), .Y(n3663) );
  AND2X1 U2951 ( .A(fifo_array[758]), .B(n5802), .Y(n966) );
  INVX1 U2952 ( .A(n966), .Y(n3664) );
  AND2X1 U2953 ( .A(fifo_array[729]), .B(n5805), .Y(n936) );
  INVX1 U2954 ( .A(n936), .Y(n3665) );
  AND2X1 U2955 ( .A(fifo_array[717]), .B(n5804), .Y(n924) );
  INVX1 U2956 ( .A(n924), .Y(n3666) );
  AND2X1 U2957 ( .A(fifo_array[689]), .B(n5807), .Y(n894) );
  INVX1 U2958 ( .A(n894), .Y(n3667) );
  AND2X1 U2959 ( .A(fifo_array[676]), .B(n5806), .Y(n881) );
  INVX1 U2960 ( .A(n881), .Y(n3668) );
  AND2X1 U2961 ( .A(fifo_array[657]), .B(n5809), .Y(n861) );
  INVX1 U2962 ( .A(n861), .Y(n3669) );
  AND2X1 U2963 ( .A(fifo_array[648]), .B(n5808), .Y(n852) );
  INVX1 U2964 ( .A(n852), .Y(n3670) );
  AND2X1 U2965 ( .A(fifo_array[635]), .B(n5808), .Y(n839) );
  INVX1 U2966 ( .A(n839), .Y(n3671) );
  AND2X1 U2967 ( .A(fifo_array[616]), .B(n5811), .Y(n819) );
  INVX1 U2968 ( .A(n819), .Y(n3672) );
  AND2X1 U2969 ( .A(fifo_array[607]), .B(n5810), .Y(n810) );
  INVX1 U2970 ( .A(n810), .Y(n3673) );
  AND2X1 U2971 ( .A(fifo_array[594]), .B(n5810), .Y(n797) );
  INVX1 U2972 ( .A(n797), .Y(n3674) );
  AND2X1 U2973 ( .A(fifo_array[575]), .B(n5813), .Y(n777) );
  INVX1 U2974 ( .A(n777), .Y(n3675) );
  AND2X1 U2975 ( .A(fifo_array[566]), .B(n5812), .Y(n768) );
  INVX1 U2976 ( .A(n768), .Y(n3676) );
  AND2X1 U2977 ( .A(fifo_array[553]), .B(n5812), .Y(n755) );
  INVX1 U2978 ( .A(n755), .Y(n3677) );
  AND2X1 U2979 ( .A(fifo_array[534]), .B(n5815), .Y(n735) );
  INVX1 U2980 ( .A(n735), .Y(n3678) );
  AND2X1 U2981 ( .A(fifo_array[528]), .B(n5814), .Y(n729) );
  INVX1 U2982 ( .A(n729), .Y(n3679) );
  AND2X1 U2983 ( .A(fifo_array[516]), .B(n5815), .Y(n717) );
  INVX1 U2984 ( .A(n717), .Y(n3680) );
  AND2X1 U2985 ( .A(fifo_array[499]), .B(n5817), .Y(n699) );
  INVX1 U2986 ( .A(n699), .Y(n3681) );
  AND2X1 U2987 ( .A(fifo_array[493]), .B(n5817), .Y(n693) );
  INVX1 U2988 ( .A(n693), .Y(n3682) );
  AND2X1 U2989 ( .A(fifo_array[458]), .B(n5819), .Y(n657) );
  INVX1 U2990 ( .A(n657), .Y(n3683) );
  AND2X1 U2991 ( .A(fifo_array[452]), .B(n5819), .Y(n651) );
  INVX1 U2992 ( .A(n651), .Y(n3684) );
  AND2X1 U2993 ( .A(fifo_array[411]), .B(n5821), .Y(n609) );
  INVX1 U2994 ( .A(n609), .Y(n3685) );
  AND2X1 U2995 ( .A(fifo_array[376]), .B(n5823), .Y(n572) );
  INVX1 U2996 ( .A(n572), .Y(n3686) );
  AND2X1 U2997 ( .A(fifo_array[370]), .B(n5823), .Y(n566) );
  INVX1 U2998 ( .A(n566), .Y(n3687) );
  AND2X1 U2999 ( .A(fifo_array[315]), .B(n5824), .Y(n509) );
  INVX1 U3000 ( .A(n509), .Y(n3688) );
  AND2X1 U3001 ( .A(fifo_array[302]), .B(n5825), .Y(n496) );
  INVX1 U3002 ( .A(n496), .Y(n3689) );
  AND2X1 U3003 ( .A(fifo_array[294]), .B(n5825), .Y(n488) );
  INVX1 U3004 ( .A(n488), .Y(n3690) );
  AND2X1 U3005 ( .A(fifo_array[277]), .B(n5826), .Y(n469) );
  INVX1 U3006 ( .A(n469), .Y(n3691) );
  AND2X1 U3007 ( .A(fifo_array[265]), .B(n5827), .Y(n457) );
  INVX1 U3008 ( .A(n457), .Y(n3692) );
  AND2X1 U3009 ( .A(fifo_array[253]), .B(n5827), .Y(n445) );
  INVX1 U3010 ( .A(n445), .Y(n3693) );
  AND2X1 U3011 ( .A(fifo_array[236]), .B(n5828), .Y(n426) );
  INVX1 U3012 ( .A(n426), .Y(n3694) );
  AND2X1 U3013 ( .A(fifo_array[224]), .B(n5829), .Y(n414) );
  INVX1 U3014 ( .A(n414), .Y(n3695) );
  AND2X1 U3015 ( .A(fifo_array[212]), .B(n5828), .Y(n402) );
  INVX1 U3016 ( .A(n402), .Y(n3696) );
  AND2X1 U3017 ( .A(fifo_array[183]), .B(n5831), .Y(n371) );
  INVX1 U3018 ( .A(n371), .Y(n3697) );
  AND2X1 U3019 ( .A(fifo_array[171]), .B(n5830), .Y(n359) );
  INVX1 U3020 ( .A(n359), .Y(n3698) );
  AND2X1 U3021 ( .A(fifo_array[143]), .B(n5833), .Y(n329) );
  INVX1 U3022 ( .A(n329), .Y(n3699) );
  AND2X1 U3023 ( .A(fifo_array[130]), .B(n5832), .Y(n316) );
  INVX1 U3024 ( .A(n316), .Y(n3700) );
  AND2X1 U3025 ( .A(fifo_array[111]), .B(n5835), .Y(n295) );
  INVX1 U3026 ( .A(n295), .Y(n3701) );
  AND2X1 U3027 ( .A(fifo_array[102]), .B(n5834), .Y(n286) );
  INVX1 U3028 ( .A(n286), .Y(n3702) );
  AND2X1 U3029 ( .A(fifo_array[89]), .B(n5834), .Y(n273) );
  INVX1 U3030 ( .A(n273), .Y(n3703) );
  AND2X1 U3031 ( .A(fifo_array[70]), .B(n5837), .Y(n252) );
  INVX1 U3032 ( .A(n252), .Y(n3704) );
  AND2X1 U3033 ( .A(fifo_array[61]), .B(n5836), .Y(n243) );
  INVX1 U3034 ( .A(n243), .Y(n3705) );
  AND2X1 U3035 ( .A(fifo_array[48]), .B(n5836), .Y(n230) );
  INVX1 U3036 ( .A(n230), .Y(n3706) );
  AND2X1 U3037 ( .A(fifo_array[29]), .B(n5839), .Y(n208) );
  INVX1 U3038 ( .A(n208), .Y(n3707) );
  AND2X1 U3039 ( .A(fifo_array[20]), .B(n5838), .Y(n199) );
  INVX1 U3040 ( .A(n199), .Y(n3708) );
  AND2X1 U3041 ( .A(fifo_array[7]), .B(n5839), .Y(n186) );
  INVX1 U3042 ( .A(n186), .Y(n3709) );
  AND2X1 U3043 ( .A(n4228), .B(n5845), .Y(n1643) );
  AND2X1 U3044 ( .A(n76), .B(n4231), .Y(n1571) );
  INVX1 U3045 ( .A(n1571), .Y(n3710) );
  AND2X1 U3046 ( .A(n5844), .B(n5773), .Y(n1589) );
  INVX1 U3047 ( .A(n1589), .Y(n3711) );
  AND2X1 U3048 ( .A(fifo_array[1317]), .B(n5776), .Y(n1539) );
  INVX1 U3049 ( .A(n1539), .Y(n3712) );
  AND2X1 U3050 ( .A(fifo_array[1305]), .B(n5777), .Y(n1527) );
  INVX1 U3051 ( .A(n1527), .Y(n3713) );
  AND2X1 U3052 ( .A(fifo_array[1286]), .B(n5779), .Y(n1507) );
  INVX1 U3053 ( .A(n1507), .Y(n3714) );
  AND2X1 U3054 ( .A(fifo_array[1274]), .B(n5778), .Y(n1495) );
  INVX1 U3055 ( .A(n1495), .Y(n3715) );
  AND2X1 U3056 ( .A(fifo_array[1262]), .B(n5779), .Y(n1483) );
  INVX1 U3057 ( .A(n1483), .Y(n3716) );
  AND2X1 U3058 ( .A(fifo_array[1245]), .B(n5780), .Y(n1465) );
  INVX1 U3059 ( .A(n1465), .Y(n3717) );
  AND2X1 U3060 ( .A(fifo_array[1236]), .B(n5781), .Y(n1456) );
  INVX1 U3061 ( .A(n1456), .Y(n3718) );
  AND2X1 U3062 ( .A(fifo_array[1223]), .B(n5781), .Y(n1443) );
  INVX1 U3063 ( .A(n1443), .Y(n3719) );
  AND2X1 U3064 ( .A(fifo_array[1193]), .B(n5782), .Y(n1412) );
  INVX1 U3065 ( .A(n1412), .Y(n3720) );
  AND2X1 U3066 ( .A(fifo_array[1180]), .B(n5783), .Y(n1399) );
  INVX1 U3067 ( .A(n1399), .Y(n3721) );
  AND2X1 U3068 ( .A(fifo_array[1163]), .B(n5784), .Y(n1381) );
  INVX1 U3069 ( .A(n1381), .Y(n3722) );
  AND2X1 U3070 ( .A(fifo_array[1154]), .B(n5785), .Y(n1372) );
  INVX1 U3071 ( .A(n1372), .Y(n3723) );
  AND2X1 U3072 ( .A(fifo_array[1141]), .B(n5785), .Y(n1359) );
  INVX1 U3073 ( .A(n1359), .Y(n3724) );
  AND2X1 U3074 ( .A(fifo_array[1120]), .B(n5786), .Y(n1337) );
  INVX1 U3075 ( .A(n1337), .Y(n3725) );
  AND2X1 U3076 ( .A(fifo_array[1111]), .B(n5787), .Y(n1328) );
  INVX1 U3077 ( .A(n1328), .Y(n3726) );
  AND2X1 U3078 ( .A(fifo_array[1098]), .B(n5787), .Y(n1315) );
  INVX1 U3079 ( .A(n1315), .Y(n3727) );
  AND2X1 U3080 ( .A(fifo_array[1089]), .B(n5789), .Y(n1305) );
  INVX1 U3081 ( .A(n1305), .Y(n3728) );
  AND2X1 U3082 ( .A(fifo_array[1073]), .B(n5788), .Y(n1289) );
  INVX1 U3083 ( .A(n1289), .Y(n3729) );
  AND2X1 U3084 ( .A(fifo_array[1061]), .B(n5788), .Y(n1277) );
  INVX1 U3085 ( .A(n1277), .Y(n3730) );
  AND2X1 U3086 ( .A(fifo_array[1046]), .B(n5791), .Y(n1260) );
  INVX1 U3087 ( .A(n1260), .Y(n3731) );
  AND2X1 U3088 ( .A(fifo_array[1040]), .B(n5791), .Y(n1254) );
  INVX1 U3089 ( .A(n1254), .Y(n3732) );
  AND2X1 U3090 ( .A(fifo_array[1003]), .B(n5792), .Y(n1216) );
  INVX1 U3091 ( .A(n1216), .Y(n3733) );
  AND2X1 U3092 ( .A(fifo_array[997]), .B(n5793), .Y(n1210) );
  INVX1 U3093 ( .A(n1210), .Y(n3734) );
  AND2X1 U3094 ( .A(fifo_array[964]), .B(n5795), .Y(n1176) );
  INVX1 U3095 ( .A(n1176), .Y(n3735) );
  AND2X1 U3096 ( .A(fifo_array[958]), .B(n5795), .Y(n1170) );
  INVX1 U3097 ( .A(n1170), .Y(n3736) );
  AND2X1 U3098 ( .A(fifo_array[915]), .B(n5797), .Y(n1126) );
  INVX1 U3099 ( .A(n1126), .Y(n3737) );
  AND2X1 U3100 ( .A(fifo_array[865]), .B(n5798), .Y(n1075) );
  INVX1 U3101 ( .A(n1075), .Y(n3738) );
  AND2X1 U3102 ( .A(fifo_array[853]), .B(n5799), .Y(n1063) );
  INVX1 U3103 ( .A(n1063), .Y(n3739) );
  AND2X1 U3104 ( .A(fifo_array[841]), .B(n5799), .Y(n1051) );
  INVX1 U3105 ( .A(n1051), .Y(n3740) );
  AND2X1 U3106 ( .A(fifo_array[819]), .B(n5800), .Y(n1028) );
  INVX1 U3107 ( .A(n1028), .Y(n3741) );
  AND2X1 U3108 ( .A(fifo_array[806]), .B(n5801), .Y(n1015) );
  INVX1 U3109 ( .A(n1015), .Y(n3742) );
  AND2X1 U3110 ( .A(fifo_array[798]), .B(n5801), .Y(n1007) );
  INVX1 U3111 ( .A(n1007), .Y(n3743) );
  AND2X1 U3112 ( .A(fifo_array[771]), .B(n5803), .Y(n979) );
  INVX1 U3113 ( .A(n979), .Y(n3744) );
  AND2X1 U3114 ( .A(fifo_array[759]), .B(n5803), .Y(n967) );
  INVX1 U3115 ( .A(n967), .Y(n3745) );
  AND2X1 U3116 ( .A(fifo_array[740]), .B(n5804), .Y(n947) );
  INVX1 U3117 ( .A(n947), .Y(n3746) );
  AND2X1 U3118 ( .A(fifo_array[728]), .B(n5805), .Y(n935) );
  INVX1 U3119 ( .A(n935), .Y(n3747) );
  AND2X1 U3120 ( .A(fifo_array[716]), .B(n5805), .Y(n923) );
  INVX1 U3121 ( .A(n923), .Y(n3748) );
  AND2X1 U3122 ( .A(fifo_array[699]), .B(n5807), .Y(n904) );
  INVX1 U3123 ( .A(n904), .Y(n3749) );
  AND2X1 U3124 ( .A(fifo_array[690]), .B(n5806), .Y(n895) );
  INVX1 U3125 ( .A(n895), .Y(n3750) );
  AND2X1 U3126 ( .A(fifo_array[677]), .B(n5807), .Y(n882) );
  INVX1 U3127 ( .A(n882), .Y(n3751) );
  AND2X1 U3128 ( .A(fifo_array[647]), .B(n5809), .Y(n851) );
  INVX1 U3129 ( .A(n851), .Y(n3752) );
  AND2X1 U3130 ( .A(fifo_array[634]), .B(n5809), .Y(n838) );
  INVX1 U3131 ( .A(n838), .Y(n3753) );
  AND2X1 U3132 ( .A(fifo_array[617]), .B(n5811), .Y(n820) );
  INVX1 U3133 ( .A(n820), .Y(n3754) );
  AND2X1 U3134 ( .A(fifo_array[608]), .B(n5810), .Y(n811) );
  INVX1 U3135 ( .A(n811), .Y(n3755) );
  AND2X1 U3136 ( .A(fifo_array[595]), .B(n5810), .Y(n798) );
  INVX1 U3137 ( .A(n798), .Y(n3756) );
  AND2X1 U3138 ( .A(fifo_array[574]), .B(n5813), .Y(n776) );
  INVX1 U3139 ( .A(n776), .Y(n3757) );
  AND2X1 U3140 ( .A(fifo_array[565]), .B(n5812), .Y(n767) );
  INVX1 U3141 ( .A(n767), .Y(n3758) );
  AND2X1 U3142 ( .A(fifo_array[552]), .B(n5812), .Y(n754) );
  INVX1 U3143 ( .A(n754), .Y(n3759) );
  AND2X1 U3144 ( .A(fifo_array[543]), .B(n5815), .Y(n744) );
  INVX1 U3145 ( .A(n744), .Y(n3760) );
  AND2X1 U3146 ( .A(fifo_array[527]), .B(n5814), .Y(n728) );
  INVX1 U3147 ( .A(n728), .Y(n3761) );
  AND2X1 U3148 ( .A(fifo_array[515]), .B(n5815), .Y(n716) );
  INVX1 U3149 ( .A(n716), .Y(n3762) );
  AND2X1 U3150 ( .A(fifo_array[500]), .B(n5816), .Y(n700) );
  INVX1 U3151 ( .A(n700), .Y(n3763) );
  AND2X1 U3152 ( .A(fifo_array[494]), .B(n5817), .Y(n694) );
  INVX1 U3153 ( .A(n694), .Y(n3764) );
  AND2X1 U3154 ( .A(fifo_array[457]), .B(n5818), .Y(n656) );
  INVX1 U3155 ( .A(n656), .Y(n3765) );
  AND2X1 U3156 ( .A(fifo_array[451]), .B(n5819), .Y(n650) );
  INVX1 U3157 ( .A(n650), .Y(n3766) );
  AND2X1 U3158 ( .A(fifo_array[418]), .B(n5821), .Y(n616) );
  INVX1 U3159 ( .A(n616), .Y(n3767) );
  AND2X1 U3160 ( .A(fifo_array[412]), .B(n5821), .Y(n610) );
  INVX1 U3161 ( .A(n610), .Y(n3768) );
  AND2X1 U3162 ( .A(fifo_array[369]), .B(n5823), .Y(n565) );
  INVX1 U3163 ( .A(n565), .Y(n3769) );
  AND2X1 U3164 ( .A(fifo_array[319]), .B(n5824), .Y(n513) );
  INVX1 U3165 ( .A(n513), .Y(n3770) );
  AND2X1 U3166 ( .A(fifo_array[307]), .B(n5825), .Y(n501) );
  INVX1 U3167 ( .A(n501), .Y(n3771) );
  AND2X1 U3168 ( .A(fifo_array[295]), .B(n5825), .Y(n489) );
  INVX1 U3169 ( .A(n489), .Y(n3772) );
  AND2X1 U3170 ( .A(fifo_array[273]), .B(n5826), .Y(n465) );
  INVX1 U3171 ( .A(n465), .Y(n3773) );
  AND2X1 U3172 ( .A(fifo_array[260]), .B(n5827), .Y(n452) );
  INVX1 U3173 ( .A(n452), .Y(n3774) );
  AND2X1 U3174 ( .A(fifo_array[252]), .B(n5827), .Y(n444) );
  INVX1 U3175 ( .A(n444), .Y(n3775) );
  AND2X1 U3176 ( .A(fifo_array[225]), .B(n5829), .Y(n415) );
  INVX1 U3177 ( .A(n415), .Y(n3776) );
  AND2X1 U3178 ( .A(fifo_array[213]), .B(n5829), .Y(n403) );
  INVX1 U3179 ( .A(n403), .Y(n3777) );
  AND2X1 U3180 ( .A(fifo_array[194]), .B(n5830), .Y(n382) );
  INVX1 U3181 ( .A(n382), .Y(n3778) );
  AND2X1 U3182 ( .A(fifo_array[182]), .B(n5831), .Y(n370) );
  INVX1 U3183 ( .A(n370), .Y(n3779) );
  AND2X1 U3184 ( .A(fifo_array[170]), .B(n5831), .Y(n358) );
  INVX1 U3185 ( .A(n358), .Y(n3780) );
  AND2X1 U3186 ( .A(fifo_array[153]), .B(n5833), .Y(n339) );
  INVX1 U3187 ( .A(n339), .Y(n3781) );
  AND2X1 U3188 ( .A(fifo_array[144]), .B(n5832), .Y(n330) );
  INVX1 U3189 ( .A(n330), .Y(n3782) );
  AND2X1 U3190 ( .A(fifo_array[131]), .B(n5833), .Y(n317) );
  INVX1 U3191 ( .A(n317), .Y(n3783) );
  AND2X1 U3192 ( .A(fifo_array[101]), .B(n5835), .Y(n285) );
  INVX1 U3193 ( .A(n285), .Y(n3784) );
  AND2X1 U3194 ( .A(fifo_array[88]), .B(n5835), .Y(n272) );
  INVX1 U3195 ( .A(n272), .Y(n3785) );
  AND2X1 U3196 ( .A(fifo_array[71]), .B(n5837), .Y(n253) );
  INVX1 U3197 ( .A(n253), .Y(n3786) );
  AND2X1 U3198 ( .A(fifo_array[62]), .B(n5836), .Y(n244) );
  INVX1 U3199 ( .A(n244), .Y(n3787) );
  AND2X1 U3200 ( .A(fifo_array[49]), .B(n5836), .Y(n231) );
  INVX1 U3201 ( .A(n231), .Y(n3788) );
  AND2X1 U3202 ( .A(fifo_array[28]), .B(n5838), .Y(n207) );
  INVX1 U3203 ( .A(n207), .Y(n3789) );
  AND2X1 U3204 ( .A(fifo_array[19]), .B(n5839), .Y(n198) );
  INVX1 U3205 ( .A(n198), .Y(n3790) );
  AND2X1 U3206 ( .A(fifo_array[6]), .B(n5839), .Y(n185) );
  INVX1 U3207 ( .A(n185), .Y(n3791) );
  AND2X1 U3208 ( .A(n77), .B(n4231), .Y(n1570) );
  INVX1 U3209 ( .A(n1570), .Y(n3792) );
  AND2X1 U3210 ( .A(n81), .B(n5773), .Y(n1588) );
  INVX1 U3211 ( .A(n1588), .Y(n3793) );
  AND2X1 U3212 ( .A(fifo_array[1323]), .B(n5777), .Y(n1545) );
  INVX1 U3213 ( .A(n1545), .Y(n3794) );
  AND2X1 U3214 ( .A(fifo_array[1310]), .B(n5776), .Y(n1532) );
  INVX1 U3215 ( .A(n1532), .Y(n3795) );
  AND2X1 U3216 ( .A(fifo_array[1302]), .B(n5777), .Y(n1524) );
  INVX1 U3217 ( .A(n1524), .Y(n3796) );
  AND2X1 U3218 ( .A(fifo_array[1285]), .B(n5779), .Y(n1506) );
  INVX1 U3219 ( .A(n1506), .Y(n3797) );
  AND2X1 U3220 ( .A(fifo_array[1273]), .B(n5778), .Y(n1494) );
  INVX1 U3221 ( .A(n1494), .Y(n3798) );
  AND2X1 U3222 ( .A(fifo_array[1261]), .B(n5779), .Y(n1482) );
  INVX1 U3223 ( .A(n1482), .Y(n3799) );
  AND2X1 U3224 ( .A(fifo_array[1246]), .B(n5780), .Y(n1466) );
  INVX1 U3225 ( .A(n1466), .Y(n3800) );
  AND2X1 U3226 ( .A(fifo_array[1237]), .B(n5781), .Y(n1457) );
  INVX1 U3227 ( .A(n1457), .Y(n3801) );
  AND2X1 U3228 ( .A(fifo_array[1224]), .B(n5781), .Y(n1444) );
  INVX1 U3229 ( .A(n1444), .Y(n3802) );
  AND2X1 U3230 ( .A(fifo_array[1205]), .B(n5782), .Y(n1424) );
  INVX1 U3231 ( .A(n1424), .Y(n3803) );
  AND2X1 U3232 ( .A(fifo_array[1196]), .B(n5783), .Y(n1415) );
  INVX1 U3233 ( .A(n1415), .Y(n3804) );
  AND2X1 U3234 ( .A(fifo_array[1183]), .B(n5783), .Y(n1402) );
  INVX1 U3235 ( .A(n1402), .Y(n3805) );
  AND2X1 U3236 ( .A(fifo_array[1151]), .B(n5784), .Y(n1369) );
  INVX1 U3237 ( .A(n1369), .Y(n3806) );
  AND2X1 U3238 ( .A(fifo_array[1138]), .B(n5785), .Y(n1356) );
  INVX1 U3239 ( .A(n1356), .Y(n3807) );
  AND2X1 U3240 ( .A(fifo_array[1119]), .B(n5786), .Y(n1336) );
  INVX1 U3241 ( .A(n1336), .Y(n3808) );
  AND2X1 U3242 ( .A(fifo_array[1110]), .B(n5787), .Y(n1327) );
  INVX1 U3243 ( .A(n1327), .Y(n3809) );
  AND2X1 U3244 ( .A(fifo_array[1097]), .B(n5787), .Y(n1314) );
  INVX1 U3245 ( .A(n1314), .Y(n3810) );
  AND2X1 U3246 ( .A(fifo_array[1086]), .B(n5789), .Y(n1302) );
  INVX1 U3247 ( .A(n1302), .Y(n3811) );
  AND2X1 U3248 ( .A(fifo_array[1072]), .B(n5789), .Y(n1288) );
  INVX1 U3249 ( .A(n1288), .Y(n3812) );
  AND2X1 U3250 ( .A(fifo_array[1060]), .B(n5789), .Y(n1276) );
  INVX1 U3251 ( .A(n1276), .Y(n3813) );
  AND2X1 U3252 ( .A(fifo_array[1041]), .B(n5790), .Y(n1255) );
  INVX1 U3253 ( .A(n1255), .Y(n3814) );
  AND2X1 U3254 ( .A(fifo_array[1006]), .B(n5793), .Y(n1219) );
  INVX1 U3255 ( .A(n1219), .Y(n3815) );
  AND2X1 U3256 ( .A(fifo_array[1000]), .B(n5793), .Y(n1213) );
  INVX1 U3257 ( .A(n1213), .Y(n3816) );
  AND2X1 U3258 ( .A(fifo_array[961]), .B(n5794), .Y(n1173) );
  INVX1 U3259 ( .A(n1173), .Y(n3817) );
  AND2X1 U3260 ( .A(fifo_array[955]), .B(n5795), .Y(n1167) );
  INVX1 U3261 ( .A(n1167), .Y(n3818) );
  AND2X1 U3262 ( .A(fifo_array[920]), .B(n5796), .Y(n1131) );
  INVX1 U3263 ( .A(n1131), .Y(n3819) );
  AND2X1 U3264 ( .A(fifo_array[914]), .B(n5797), .Y(n1125) );
  INVX1 U3265 ( .A(n1125), .Y(n3820) );
  AND2X1 U3266 ( .A(fifo_array[866]), .B(n5798), .Y(n1076) );
  INVX1 U3267 ( .A(n1076), .Y(n3821) );
  AND2X1 U3268 ( .A(fifo_array[854]), .B(n5799), .Y(n1064) );
  INVX1 U3269 ( .A(n1064), .Y(n3822) );
  AND2X1 U3270 ( .A(fifo_array[842]), .B(n5798), .Y(n1052) );
  INVX1 U3271 ( .A(n1052), .Y(n3823) );
  AND2X1 U3272 ( .A(fifo_array[813]), .B(n5801), .Y(n1022) );
  INVX1 U3273 ( .A(n1022), .Y(n3824) );
  AND2X1 U3274 ( .A(fifo_array[801]), .B(n5800), .Y(n1010) );
  INVX1 U3275 ( .A(n1010), .Y(n3825) );
  AND2X1 U3276 ( .A(fifo_array[777]), .B(n5802), .Y(n985) );
  INVX1 U3277 ( .A(n985), .Y(n3826) );
  AND2X1 U3278 ( .A(fifo_array[764]), .B(n5803), .Y(n972) );
  INVX1 U3279 ( .A(n972), .Y(n3827) );
  AND2X1 U3280 ( .A(fifo_array[756]), .B(n5803), .Y(n964) );
  INVX1 U3281 ( .A(n964), .Y(n3828) );
  AND2X1 U3282 ( .A(fifo_array[739]), .B(n5804), .Y(n946) );
  INVX1 U3283 ( .A(n946), .Y(n3829) );
  AND2X1 U3284 ( .A(fifo_array[727]), .B(n5805), .Y(n934) );
  INVX1 U3285 ( .A(n934), .Y(n3830) );
  AND2X1 U3286 ( .A(fifo_array[715]), .B(n5805), .Y(n922) );
  INVX1 U3287 ( .A(n922), .Y(n3831) );
  AND2X1 U3288 ( .A(fifo_array[700]), .B(n5807), .Y(n905) );
  INVX1 U3289 ( .A(n905), .Y(n3832) );
  AND2X1 U3290 ( .A(fifo_array[691]), .B(n5806), .Y(n896) );
  INVX1 U3291 ( .A(n896), .Y(n3833) );
  AND2X1 U3292 ( .A(fifo_array[678]), .B(n5806), .Y(n883) );
  INVX1 U3293 ( .A(n883), .Y(n3834) );
  AND2X1 U3294 ( .A(fifo_array[659]), .B(n5809), .Y(n863) );
  INVX1 U3295 ( .A(n863), .Y(n3835) );
  AND2X1 U3296 ( .A(fifo_array[650]), .B(n5808), .Y(n854) );
  INVX1 U3297 ( .A(n854), .Y(n3836) );
  AND2X1 U3298 ( .A(fifo_array[637]), .B(n5808), .Y(n841) );
  INVX1 U3299 ( .A(n841), .Y(n3837) );
  AND2X1 U3300 ( .A(fifo_array[605]), .B(n5811), .Y(n808) );
  INVX1 U3301 ( .A(n808), .Y(n3838) );
  AND2X1 U3302 ( .A(fifo_array[592]), .B(n5810), .Y(n795) );
  INVX1 U3303 ( .A(n795), .Y(n3839) );
  AND2X1 U3304 ( .A(fifo_array[573]), .B(n5813), .Y(n775) );
  INVX1 U3305 ( .A(n775), .Y(n3840) );
  AND2X1 U3306 ( .A(fifo_array[564]), .B(n5812), .Y(n766) );
  INVX1 U3307 ( .A(n766), .Y(n3841) );
  AND2X1 U3308 ( .A(fifo_array[551]), .B(n5812), .Y(n753) );
  INVX1 U3309 ( .A(n753), .Y(n3842) );
  AND2X1 U3310 ( .A(fifo_array[540]), .B(n5814), .Y(n741) );
  INVX1 U3311 ( .A(n741), .Y(n3843) );
  AND2X1 U3312 ( .A(fifo_array[526]), .B(n5814), .Y(n727) );
  INVX1 U3313 ( .A(n727), .Y(n3844) );
  AND2X1 U3314 ( .A(fifo_array[514]), .B(n5815), .Y(n715) );
  INVX1 U3315 ( .A(n715), .Y(n3845) );
  AND2X1 U3316 ( .A(fifo_array[495]), .B(n5817), .Y(n695) );
  INVX1 U3317 ( .A(n695), .Y(n3846) );
  AND2X1 U3318 ( .A(fifo_array[460]), .B(n5819), .Y(n659) );
  INVX1 U3319 ( .A(n659), .Y(n3847) );
  AND2X1 U3320 ( .A(fifo_array[454]), .B(n5819), .Y(n653) );
  INVX1 U3321 ( .A(n653), .Y(n3848) );
  AND2X1 U3322 ( .A(fifo_array[415]), .B(n5820), .Y(n613) );
  INVX1 U3323 ( .A(n613), .Y(n3849) );
  AND2X1 U3324 ( .A(fifo_array[409]), .B(n5821), .Y(n607) );
  INVX1 U3325 ( .A(n607), .Y(n3850) );
  AND2X1 U3326 ( .A(fifo_array[374]), .B(n5822), .Y(n570) );
  INVX1 U3327 ( .A(n570), .Y(n3851) );
  AND2X1 U3328 ( .A(fifo_array[368]), .B(n5823), .Y(n564) );
  INVX1 U3329 ( .A(n564), .Y(n3852) );
  AND2X1 U3330 ( .A(fifo_array[320]), .B(n5824), .Y(n514) );
  INVX1 U3331 ( .A(n514), .Y(n3853) );
  AND2X1 U3332 ( .A(fifo_array[308]), .B(n5825), .Y(n502) );
  INVX1 U3333 ( .A(n502), .Y(n3854) );
  AND2X1 U3334 ( .A(fifo_array[296]), .B(n5824), .Y(n490) );
  INVX1 U3335 ( .A(n490), .Y(n3855) );
  AND2X1 U3336 ( .A(fifo_array[267]), .B(n5827), .Y(n459) );
  INVX1 U3337 ( .A(n459), .Y(n3856) );
  AND2X1 U3338 ( .A(fifo_array[255]), .B(n5826), .Y(n447) );
  INVX1 U3339 ( .A(n447), .Y(n3857) );
  AND2X1 U3340 ( .A(fifo_array[231]), .B(n5828), .Y(n421) );
  INVX1 U3341 ( .A(n421), .Y(n3858) );
  AND2X1 U3342 ( .A(fifo_array[218]), .B(n5829), .Y(n408) );
  INVX1 U3343 ( .A(n408), .Y(n3859) );
  AND2X1 U3344 ( .A(fifo_array[210]), .B(n5829), .Y(n400) );
  INVX1 U3345 ( .A(n400), .Y(n3860) );
  AND2X1 U3346 ( .A(fifo_array[193]), .B(n5830), .Y(n381) );
  INVX1 U3347 ( .A(n381), .Y(n3861) );
  AND2X1 U3348 ( .A(fifo_array[181]), .B(n5831), .Y(n369) );
  INVX1 U3349 ( .A(n369), .Y(n3862) );
  AND2X1 U3350 ( .A(fifo_array[169]), .B(n5831), .Y(n357) );
  INVX1 U3351 ( .A(n357), .Y(n3863) );
  AND2X1 U3352 ( .A(fifo_array[154]), .B(n5833), .Y(n340) );
  INVX1 U3353 ( .A(n340), .Y(n3864) );
  AND2X1 U3354 ( .A(fifo_array[145]), .B(n5832), .Y(n331) );
  INVX1 U3355 ( .A(n331), .Y(n3865) );
  AND2X1 U3356 ( .A(fifo_array[132]), .B(n5832), .Y(n318) );
  INVX1 U3357 ( .A(n318), .Y(n3866) );
  AND2X1 U3358 ( .A(fifo_array[113]), .B(n5835), .Y(n297) );
  INVX1 U3359 ( .A(n297), .Y(n3867) );
  AND2X1 U3360 ( .A(fifo_array[104]), .B(n5834), .Y(n288) );
  INVX1 U3361 ( .A(n288), .Y(n3868) );
  AND2X1 U3362 ( .A(fifo_array[91]), .B(n5834), .Y(n275) );
  INVX1 U3363 ( .A(n275), .Y(n3869) );
  AND2X1 U3364 ( .A(fifo_array[59]), .B(n5837), .Y(n241) );
  INVX1 U3365 ( .A(n241), .Y(n3870) );
  AND2X1 U3366 ( .A(fifo_array[46]), .B(n5836), .Y(n228) );
  INVX1 U3367 ( .A(n228), .Y(n3871) );
  AND2X1 U3368 ( .A(fifo_array[27]), .B(n5838), .Y(n206) );
  INVX1 U3369 ( .A(n206), .Y(n3872) );
  AND2X1 U3370 ( .A(fifo_array[18]), .B(n5839), .Y(n197) );
  INVX1 U3371 ( .A(n197), .Y(n3873) );
  AND2X1 U3372 ( .A(fifo_array[5]), .B(n5839), .Y(n184) );
  INVX1 U3373 ( .A(n184), .Y(n3874) );
  AND2X1 U3374 ( .A(n5845), .B(n4321), .Y(n1636) );
  INVX1 U3375 ( .A(n1636), .Y(n3875) );
  AND2X1 U3376 ( .A(n78), .B(n4231), .Y(n1569) );
  INVX1 U3377 ( .A(n1569), .Y(n3876) );
  AND2X1 U3378 ( .A(n82), .B(n5775), .Y(n1587) );
  INVX1 U3379 ( .A(n1587), .Y(n3877) );
  AND2X1 U3380 ( .A(fifo_array[1327]), .B(n5777), .Y(n1549) );
  INVX1 U3381 ( .A(n1549), .Y(n3878) );
  AND2X1 U3382 ( .A(fifo_array[1315]), .B(n5776), .Y(n1537) );
  INVX1 U3383 ( .A(n1537), .Y(n3879) );
  AND2X1 U3384 ( .A(fifo_array[1303]), .B(n5777), .Y(n1525) );
  INVX1 U3385 ( .A(n1525), .Y(n3880) );
  AND2X1 U3386 ( .A(fifo_array[1281]), .B(n5779), .Y(n1502) );
  INVX1 U3387 ( .A(n1502), .Y(n3881) );
  AND2X1 U3388 ( .A(fifo_array[1268]), .B(n5778), .Y(n1489) );
  INVX1 U3389 ( .A(n1489), .Y(n3882) );
  AND2X1 U3390 ( .A(fifo_array[1260]), .B(n5779), .Y(n1481) );
  INVX1 U3391 ( .A(n1481), .Y(n3883) );
  AND2X1 U3392 ( .A(fifo_array[1247]), .B(n5780), .Y(n1467) );
  INVX1 U3393 ( .A(n1467), .Y(n3884) );
  AND2X1 U3394 ( .A(fifo_array[1238]), .B(n5781), .Y(n1458) );
  INVX1 U3395 ( .A(n1458), .Y(n3885) );
  AND2X1 U3396 ( .A(fifo_array[1225]), .B(n5781), .Y(n1445) );
  INVX1 U3397 ( .A(n1445), .Y(n3886) );
  AND2X1 U3398 ( .A(fifo_array[1204]), .B(n5782), .Y(n1423) );
  INVX1 U3399 ( .A(n1423), .Y(n3887) );
  AND2X1 U3400 ( .A(fifo_array[1195]), .B(n5783), .Y(n1414) );
  INVX1 U3401 ( .A(n1414), .Y(n3888) );
  AND2X1 U3402 ( .A(fifo_array[1182]), .B(n5783), .Y(n1401) );
  INVX1 U3403 ( .A(n1401), .Y(n3889) );
  AND2X1 U3404 ( .A(fifo_array[1161]), .B(n5784), .Y(n1379) );
  INVX1 U3405 ( .A(n1379), .Y(n3890) );
  AND2X1 U3406 ( .A(fifo_array[1152]), .B(n5785), .Y(n1370) );
  INVX1 U3407 ( .A(n1370), .Y(n3891) );
  AND2X1 U3408 ( .A(fifo_array[1139]), .B(n5785), .Y(n1357) );
  INVX1 U3409 ( .A(n1357), .Y(n3892) );
  AND2X1 U3410 ( .A(fifo_array[1109]), .B(n5786), .Y(n1326) );
  INVX1 U3411 ( .A(n1326), .Y(n3893) );
  AND2X1 U3412 ( .A(fifo_array[1096]), .B(n5787), .Y(n1313) );
  INVX1 U3413 ( .A(n1313), .Y(n3894) );
  AND2X1 U3414 ( .A(fifo_array[1066]), .B(n5789), .Y(n1282) );
  INVX1 U3415 ( .A(n1282), .Y(n3895) );
  AND2X1 U3416 ( .A(fifo_array[1059]), .B(n5788), .Y(n1275) );
  INVX1 U3417 ( .A(n1275), .Y(n3896) );
  AND2X1 U3418 ( .A(fifo_array[1048]), .B(n5791), .Y(n1262) );
  INVX1 U3419 ( .A(n1262), .Y(n3897) );
  AND2X1 U3420 ( .A(fifo_array[1042]), .B(n5791), .Y(n1256) );
  INVX1 U3421 ( .A(n1256), .Y(n3898) );
  AND2X1 U3422 ( .A(fifo_array[999]), .B(n5793), .Y(n1212) );
  INVX1 U3423 ( .A(n1212), .Y(n3899) );
  AND2X1 U3424 ( .A(fifo_array[962]), .B(n5795), .Y(n1174) );
  INVX1 U3425 ( .A(n1174), .Y(n3900) );
  AND2X1 U3426 ( .A(fifo_array[956]), .B(n5795), .Y(n1168) );
  INVX1 U3427 ( .A(n1168), .Y(n3901) );
  AND2X1 U3428 ( .A(fifo_array[919]), .B(n5797), .Y(n1130) );
  INVX1 U3429 ( .A(n1130), .Y(n3902) );
  AND2X1 U3430 ( .A(fifo_array[913]), .B(n5797), .Y(n1124) );
  INVX1 U3431 ( .A(n1124), .Y(n3903) );
  AND2X1 U3432 ( .A(fifo_array[855]), .B(n5799), .Y(n1065) );
  INVX1 U3433 ( .A(n1065), .Y(n3904) );
  AND2X1 U3434 ( .A(fifo_array[843]), .B(n5799), .Y(n1053) );
  INVX1 U3435 ( .A(n1053), .Y(n3905) );
  AND2X1 U3436 ( .A(fifo_array[824]), .B(n5800), .Y(n1033) );
  INVX1 U3437 ( .A(n1033), .Y(n3906) );
  AND2X1 U3438 ( .A(fifo_array[812]), .B(n5801), .Y(n1021) );
  INVX1 U3439 ( .A(n1021), .Y(n3907) );
  AND2X1 U3440 ( .A(fifo_array[800]), .B(n5801), .Y(n1009) );
  INVX1 U3441 ( .A(n1009), .Y(n3908) );
  AND2X1 U3442 ( .A(fifo_array[781]), .B(n5802), .Y(n989) );
  INVX1 U3443 ( .A(n989), .Y(n3909) );
  AND2X1 U3444 ( .A(fifo_array[769]), .B(n5803), .Y(n977) );
  INVX1 U3445 ( .A(n977), .Y(n3910) );
  AND2X1 U3446 ( .A(fifo_array[757]), .B(n5803), .Y(n965) );
  INVX1 U3447 ( .A(n965), .Y(n3911) );
  AND2X1 U3448 ( .A(fifo_array[735]), .B(n5804), .Y(n942) );
  INVX1 U3449 ( .A(n942), .Y(n3912) );
  AND2X1 U3450 ( .A(fifo_array[722]), .B(n5805), .Y(n929) );
  INVX1 U3451 ( .A(n929), .Y(n3913) );
  AND2X1 U3452 ( .A(fifo_array[714]), .B(n5805), .Y(n921) );
  INVX1 U3453 ( .A(n921), .Y(n3914) );
  AND2X1 U3454 ( .A(fifo_array[701]), .B(n5807), .Y(n906) );
  INVX1 U3455 ( .A(n906), .Y(n3915) );
  AND2X1 U3456 ( .A(fifo_array[692]), .B(n5806), .Y(n897) );
  INVX1 U3457 ( .A(n897), .Y(n3916) );
  AND2X1 U3458 ( .A(fifo_array[679]), .B(n5806), .Y(n884) );
  INVX1 U3459 ( .A(n884), .Y(n3917) );
  AND2X1 U3460 ( .A(fifo_array[658]), .B(n5809), .Y(n862) );
  INVX1 U3461 ( .A(n862), .Y(n3918) );
  AND2X1 U3462 ( .A(fifo_array[649]), .B(n5808), .Y(n853) );
  INVX1 U3463 ( .A(n853), .Y(n3919) );
  AND2X1 U3464 ( .A(fifo_array[636]), .B(n5808), .Y(n840) );
  INVX1 U3465 ( .A(n840), .Y(n3920) );
  AND2X1 U3466 ( .A(fifo_array[615]), .B(n5811), .Y(n818) );
  INVX1 U3467 ( .A(n818), .Y(n3921) );
  AND2X1 U3468 ( .A(fifo_array[606]), .B(n5810), .Y(n809) );
  INVX1 U3469 ( .A(n809), .Y(n3922) );
  AND2X1 U3470 ( .A(fifo_array[593]), .B(n5811), .Y(n796) );
  INVX1 U3471 ( .A(n796), .Y(n3923) );
  AND2X1 U3472 ( .A(fifo_array[563]), .B(n5813), .Y(n765) );
  INVX1 U3473 ( .A(n765), .Y(n3924) );
  AND2X1 U3474 ( .A(fifo_array[550]), .B(n5813), .Y(n752) );
  INVX1 U3475 ( .A(n752), .Y(n3925) );
  AND2X1 U3476 ( .A(fifo_array[520]), .B(n5815), .Y(n721) );
  INVX1 U3477 ( .A(n721), .Y(n3926) );
  AND2X1 U3478 ( .A(fifo_array[513]), .B(n5815), .Y(n714) );
  INVX1 U3479 ( .A(n714), .Y(n3927) );
  AND2X1 U3480 ( .A(fifo_array[502]), .B(n5817), .Y(n702) );
  INVX1 U3481 ( .A(n702), .Y(n3928) );
  AND2X1 U3482 ( .A(fifo_array[496]), .B(n5817), .Y(n696) );
  INVX1 U3483 ( .A(n696), .Y(n3929) );
  AND2X1 U3484 ( .A(fifo_array[453]), .B(n5819), .Y(n652) );
  INVX1 U3485 ( .A(n652), .Y(n3930) );
  AND2X1 U3486 ( .A(fifo_array[416]), .B(n5821), .Y(n614) );
  INVX1 U3487 ( .A(n614), .Y(n3931) );
  AND2X1 U3488 ( .A(fifo_array[410]), .B(n5821), .Y(n608) );
  INVX1 U3489 ( .A(n608), .Y(n3932) );
  AND2X1 U3490 ( .A(fifo_array[373]), .B(n5823), .Y(n569) );
  INVX1 U3491 ( .A(n569), .Y(n3933) );
  AND2X1 U3492 ( .A(fifo_array[367]), .B(n5823), .Y(n563) );
  INVX1 U3493 ( .A(n563), .Y(n3934) );
  AND2X1 U3494 ( .A(fifo_array[309]), .B(n5825), .Y(n503) );
  INVX1 U3495 ( .A(n503), .Y(n3935) );
  AND2X1 U3496 ( .A(fifo_array[297]), .B(n5825), .Y(n491) );
  INVX1 U3497 ( .A(n491), .Y(n3936) );
  AND2X1 U3498 ( .A(fifo_array[278]), .B(n5826), .Y(n470) );
  INVX1 U3499 ( .A(n470), .Y(n3937) );
  AND2X1 U3500 ( .A(fifo_array[266]), .B(n5827), .Y(n458) );
  INVX1 U3501 ( .A(n458), .Y(n3938) );
  AND2X1 U3502 ( .A(fifo_array[254]), .B(n5827), .Y(n446) );
  INVX1 U3503 ( .A(n446), .Y(n3939) );
  AND2X1 U3504 ( .A(fifo_array[235]), .B(n5828), .Y(n425) );
  INVX1 U3505 ( .A(n425), .Y(n3940) );
  AND2X1 U3506 ( .A(fifo_array[223]), .B(n5829), .Y(n413) );
  INVX1 U3507 ( .A(n413), .Y(n3941) );
  AND2X1 U3508 ( .A(fifo_array[211]), .B(n5829), .Y(n401) );
  INVX1 U3509 ( .A(n401), .Y(n3942) );
  AND2X1 U3510 ( .A(fifo_array[189]), .B(n5830), .Y(n377) );
  INVX1 U3511 ( .A(n377), .Y(n3943) );
  AND2X1 U3512 ( .A(fifo_array[176]), .B(n5831), .Y(n364) );
  INVX1 U3513 ( .A(n364), .Y(n3944) );
  AND2X1 U3514 ( .A(fifo_array[168]), .B(n5831), .Y(n356) );
  INVX1 U3515 ( .A(n356), .Y(n3945) );
  AND2X1 U3516 ( .A(fifo_array[155]), .B(n5833), .Y(n341) );
  INVX1 U3517 ( .A(n341), .Y(n3946) );
  AND2X1 U3518 ( .A(fifo_array[146]), .B(n5832), .Y(n332) );
  INVX1 U3519 ( .A(n332), .Y(n3947) );
  AND2X1 U3520 ( .A(fifo_array[133]), .B(n5832), .Y(n319) );
  INVX1 U3521 ( .A(n319), .Y(n3948) );
  AND2X1 U3522 ( .A(fifo_array[112]), .B(n5835), .Y(n296) );
  INVX1 U3523 ( .A(n296), .Y(n3949) );
  AND2X1 U3524 ( .A(fifo_array[103]), .B(n5834), .Y(n287) );
  INVX1 U3525 ( .A(n287), .Y(n3950) );
  AND2X1 U3526 ( .A(fifo_array[90]), .B(n5834), .Y(n274) );
  INVX1 U3527 ( .A(n274), .Y(n3951) );
  AND2X1 U3528 ( .A(fifo_array[69]), .B(n5837), .Y(n251) );
  INVX1 U3529 ( .A(n251), .Y(n3952) );
  AND2X1 U3530 ( .A(fifo_array[60]), .B(n5836), .Y(n242) );
  INVX1 U3531 ( .A(n242), .Y(n3953) );
  AND2X1 U3532 ( .A(fifo_array[47]), .B(n5837), .Y(n229) );
  INVX1 U3533 ( .A(n229), .Y(n3954) );
  AND2X1 U3534 ( .A(fifo_array[17]), .B(n5839), .Y(n196) );
  INVX1 U3535 ( .A(n196), .Y(n3955) );
  AND2X1 U3536 ( .A(fifo_array[4]), .B(n5839), .Y(n183) );
  INVX1 U3537 ( .A(n183), .Y(n3956) );
  BUFX2 U3538 ( .A(n1633), .Y(n3957) );
  INVX1 U3539 ( .A(n1645), .Y(n3958) );
  BUFX2 U3540 ( .A(n1644), .Y(n3959) );
  BUFX2 U3541 ( .A(n1646), .Y(n3960) );
  AND2X1 U3542 ( .A(n79), .B(n4231), .Y(n1567) );
  INVX1 U3543 ( .A(n1567), .Y(n3961) );
  AND2X1 U3544 ( .A(n83), .B(n5773), .Y(n1586) );
  INVX1 U3545 ( .A(n1586), .Y(n3962) );
  AND2X1 U3546 ( .A(fifo_array[1330]), .B(n5776), .Y(n1552) );
  INVX1 U3547 ( .A(n1552), .Y(n3963) );
  AND2X1 U3548 ( .A(fifo_array[1321]), .B(n5776), .Y(n1543) );
  INVX1 U3549 ( .A(n1543), .Y(n3964) );
  AND2X1 U3550 ( .A(fifo_array[1308]), .B(n5777), .Y(n1530) );
  INVX1 U3551 ( .A(n1530), .Y(n3965) );
  AND2X1 U3552 ( .A(fifo_array[1289]), .B(n5778), .Y(n1510) );
  INVX1 U3553 ( .A(n1510), .Y(n3966) );
  AND2X1 U3554 ( .A(fifo_array[1280]), .B(n5778), .Y(n1501) );
  INVX1 U3555 ( .A(n1501), .Y(n3967) );
  AND2X1 U3556 ( .A(fifo_array[1267]), .B(n5779), .Y(n1488) );
  INVX1 U3557 ( .A(n1488), .Y(n3968) );
  AND2X1 U3558 ( .A(fifo_array[1239]), .B(n5780), .Y(n1459) );
  INVX1 U3559 ( .A(n1459), .Y(n3969) );
  AND2X1 U3560 ( .A(fifo_array[1226]), .B(n5780), .Y(n1446) );
  INVX1 U3561 ( .A(n1446), .Y(n3970) );
  AND2X1 U3562 ( .A(fifo_array[1218]), .B(n5781), .Y(n1438) );
  INVX1 U3563 ( .A(n1438), .Y(n3971) );
  AND2X1 U3564 ( .A(fifo_array[1201]), .B(n5782), .Y(n1420) );
  INVX1 U3565 ( .A(n1420), .Y(n3972) );
  AND2X1 U3566 ( .A(fifo_array[1189]), .B(n5782), .Y(n1408) );
  INVX1 U3567 ( .A(n1408), .Y(n3973) );
  AND2X1 U3568 ( .A(fifo_array[1177]), .B(n5783), .Y(n1396) );
  INVX1 U3569 ( .A(n1396), .Y(n3974) );
  AND2X1 U3570 ( .A(fifo_array[1160]), .B(n5784), .Y(n1378) );
  INVX1 U3571 ( .A(n1378), .Y(n3975) );
  AND2X1 U3572 ( .A(fifo_array[1148]), .B(n5784), .Y(n1366) );
  INVX1 U3573 ( .A(n1366), .Y(n3976) );
  AND2X1 U3574 ( .A(fifo_array[1136]), .B(n5785), .Y(n1354) );
  INVX1 U3575 ( .A(n1354), .Y(n3977) );
  AND2X1 U3576 ( .A(fifo_array[1107]), .B(n5786), .Y(n1324) );
  INVX1 U3577 ( .A(n1324), .Y(n3978) );
  AND2X1 U3578 ( .A(fifo_array[1095]), .B(n5787), .Y(n1312) );
  INVX1 U3579 ( .A(n1312), .Y(n3979) );
  AND2X1 U3580 ( .A(fifo_array[1090]), .B(n5789), .Y(n1306) );
  INVX1 U3581 ( .A(n1306), .Y(n3980) );
  AND2X1 U3582 ( .A(fifo_array[1084]), .B(n5789), .Y(n1300) );
  INVX1 U3583 ( .A(n1300), .Y(n3981) );
  AND2X1 U3584 ( .A(fifo_array[1024]), .B(n5791), .Y(n1238) );
  INVX1 U3585 ( .A(n1238), .Y(n3982) );
  AND2X1 U3586 ( .A(fifo_array[1017]), .B(n5790), .Y(n1231) );
  INVX1 U3587 ( .A(n1231), .Y(n3983) );
  AND2X1 U3588 ( .A(fifo_array[1002]), .B(n5792), .Y(n1215) );
  INVX1 U3589 ( .A(n1215), .Y(n3984) );
  AND2X1 U3590 ( .A(fifo_array[988]), .B(n5792), .Y(n1201) );
  INVX1 U3591 ( .A(n1201), .Y(n3985) );
  AND2X1 U3592 ( .A(fifo_array[976]), .B(n5793), .Y(n1189) );
  INVX1 U3593 ( .A(n1189), .Y(n3986) );
  AND2X1 U3594 ( .A(fifo_array[963]), .B(n5794), .Y(n1175) );
  INVX1 U3595 ( .A(n1175), .Y(n3987) );
  AND2X1 U3596 ( .A(fifo_array[947]), .B(n5794), .Y(n1159) );
  INVX1 U3597 ( .A(n1159), .Y(n3988) );
  AND2X1 U3598 ( .A(fifo_array[935]), .B(n5795), .Y(n1147) );
  INVX1 U3599 ( .A(n1147), .Y(n3989) );
  AND2X1 U3600 ( .A(fifo_array[912]), .B(n5797), .Y(n1123) );
  INVX1 U3601 ( .A(n1123), .Y(n3990) );
  AND2X1 U3602 ( .A(fifo_array[906]), .B(n5796), .Y(n1117) );
  INVX1 U3603 ( .A(n1117), .Y(n3991) );
  AND2X1 U3604 ( .A(fifo_array[894]), .B(n5797), .Y(n1105) );
  INVX1 U3605 ( .A(n1105), .Y(n3992) );
  AND2X1 U3606 ( .A(fifo_array[857]), .B(n5799), .Y(n1067) );
  INVX1 U3607 ( .A(n1067), .Y(n3993) );
  AND2X1 U3608 ( .A(fifo_array[844]), .B(n5798), .Y(n1054) );
  INVX1 U3609 ( .A(n1054), .Y(n3994) );
  AND2X1 U3610 ( .A(fifo_array[825]), .B(n5801), .Y(n1034) );
  INVX1 U3611 ( .A(n1034), .Y(n3995) );
  AND2X1 U3612 ( .A(fifo_array[816]), .B(n5800), .Y(n1025) );
  INVX1 U3613 ( .A(n1025), .Y(n3996) );
  AND2X1 U3614 ( .A(fifo_array[803]), .B(n5800), .Y(n1012) );
  INVX1 U3615 ( .A(n1012), .Y(n3997) );
  AND2X1 U3616 ( .A(fifo_array[784]), .B(n5803), .Y(n992) );
  INVX1 U3617 ( .A(n992), .Y(n3998) );
  AND2X1 U3618 ( .A(fifo_array[775]), .B(n5802), .Y(n983) );
  INVX1 U3619 ( .A(n983), .Y(n3999) );
  AND2X1 U3620 ( .A(fifo_array[762]), .B(n5802), .Y(n970) );
  INVX1 U3621 ( .A(n970), .Y(n4000) );
  AND2X1 U3622 ( .A(fifo_array[743]), .B(n5805), .Y(n950) );
  INVX1 U3623 ( .A(n950), .Y(n4001) );
  AND2X1 U3624 ( .A(fifo_array[734]), .B(n5804), .Y(n941) );
  INVX1 U3625 ( .A(n941), .Y(n4002) );
  AND2X1 U3626 ( .A(fifo_array[721]), .B(n5804), .Y(n928) );
  INVX1 U3627 ( .A(n928), .Y(n4003) );
  AND2X1 U3628 ( .A(fifo_array[693]), .B(n5806), .Y(n898) );
  INVX1 U3629 ( .A(n898), .Y(n4004) );
  AND2X1 U3630 ( .A(fifo_array[680]), .B(n5807), .Y(n885) );
  INVX1 U3631 ( .A(n885), .Y(n4005) );
  AND2X1 U3632 ( .A(fifo_array[672]), .B(n5807), .Y(n877) );
  INVX1 U3633 ( .A(n877), .Y(n4006) );
  AND2X1 U3634 ( .A(fifo_array[655]), .B(n5808), .Y(n859) );
  INVX1 U3635 ( .A(n859), .Y(n4007) );
  AND2X1 U3636 ( .A(fifo_array[643]), .B(n5809), .Y(n847) );
  INVX1 U3637 ( .A(n847), .Y(n4008) );
  AND2X1 U3638 ( .A(fifo_array[631]), .B(n5809), .Y(n835) );
  INVX1 U3639 ( .A(n835), .Y(n4009) );
  AND2X1 U3640 ( .A(fifo_array[614]), .B(n5810), .Y(n817) );
  INVX1 U3641 ( .A(n817), .Y(n4010) );
  AND2X1 U3642 ( .A(fifo_array[602]), .B(n5811), .Y(n805) );
  INVX1 U3643 ( .A(n805), .Y(n4011) );
  AND2X1 U3644 ( .A(fifo_array[590]), .B(n5810), .Y(n793) );
  INVX1 U3645 ( .A(n793), .Y(n4012) );
  AND2X1 U3646 ( .A(fifo_array[561]), .B(n5813), .Y(n763) );
  INVX1 U3647 ( .A(n763), .Y(n4013) );
  AND2X1 U3648 ( .A(fifo_array[549]), .B(n5812), .Y(n751) );
  INVX1 U3649 ( .A(n751), .Y(n4014) );
  AND2X1 U3650 ( .A(fifo_array[544]), .B(n5814), .Y(n745) );
  INVX1 U3651 ( .A(n745), .Y(n4015) );
  AND2X1 U3652 ( .A(fifo_array[538]), .B(n5815), .Y(n739) );
  INVX1 U3653 ( .A(n739), .Y(n4016) );
  AND2X1 U3654 ( .A(fifo_array[478]), .B(n5816), .Y(n678) );
  INVX1 U3655 ( .A(n678), .Y(n4017) );
  AND2X1 U3656 ( .A(fifo_array[471]), .B(n5817), .Y(n671) );
  INVX1 U3657 ( .A(n671), .Y(n4018) );
  AND2X1 U3658 ( .A(fifo_array[456]), .B(n5818), .Y(n655) );
  INVX1 U3659 ( .A(n655), .Y(n4019) );
  AND2X1 U3660 ( .A(fifo_array[442]), .B(n5818), .Y(n641) );
  INVX1 U3661 ( .A(n641), .Y(n4020) );
  AND2X1 U3662 ( .A(fifo_array[430]), .B(n5819), .Y(n629) );
  INVX1 U3663 ( .A(n629), .Y(n4021) );
  AND2X1 U3664 ( .A(fifo_array[417]), .B(n5820), .Y(n615) );
  INVX1 U3665 ( .A(n615), .Y(n4022) );
  AND2X1 U3666 ( .A(fifo_array[401]), .B(n5820), .Y(n599) );
  INVX1 U3667 ( .A(n599), .Y(n4023) );
  AND2X1 U3668 ( .A(fifo_array[389]), .B(n5821), .Y(n587) );
  INVX1 U3669 ( .A(n587), .Y(n4024) );
  AND2X1 U3670 ( .A(fifo_array[366]), .B(n5823), .Y(n562) );
  INVX1 U3671 ( .A(n562), .Y(n4025) );
  AND2X1 U3672 ( .A(fifo_array[360]), .B(n5822), .Y(n556) );
  INVX1 U3673 ( .A(n556), .Y(n4026) );
  AND2X1 U3674 ( .A(fifo_array[348]), .B(n5823), .Y(n544) );
  INVX1 U3675 ( .A(n544), .Y(n4027) );
  AND2X1 U3676 ( .A(fifo_array[311]), .B(n5825), .Y(n505) );
  INVX1 U3677 ( .A(n505), .Y(n4028) );
  AND2X1 U3678 ( .A(fifo_array[298]), .B(n5824), .Y(n492) );
  INVX1 U3679 ( .A(n492), .Y(n4029) );
  AND2X1 U3680 ( .A(fifo_array[279]), .B(n5827), .Y(n471) );
  INVX1 U3681 ( .A(n471), .Y(n4030) );
  AND2X1 U3682 ( .A(fifo_array[270]), .B(n5826), .Y(n462) );
  INVX1 U3683 ( .A(n462), .Y(n4031) );
  AND2X1 U3684 ( .A(fifo_array[257]), .B(n5826), .Y(n449) );
  INVX1 U3685 ( .A(n449), .Y(n4032) );
  AND2X1 U3686 ( .A(fifo_array[238]), .B(n5829), .Y(n428) );
  INVX1 U3687 ( .A(n428), .Y(n4033) );
  AND2X1 U3688 ( .A(fifo_array[229]), .B(n5828), .Y(n419) );
  INVX1 U3689 ( .A(n419), .Y(n4034) );
  AND2X1 U3690 ( .A(fifo_array[216]), .B(n5828), .Y(n406) );
  INVX1 U3691 ( .A(n406), .Y(n4035) );
  AND2X1 U3692 ( .A(fifo_array[197]), .B(n5831), .Y(n385) );
  INVX1 U3693 ( .A(n385), .Y(n4036) );
  AND2X1 U3694 ( .A(fifo_array[188]), .B(n5830), .Y(n376) );
  INVX1 U3695 ( .A(n376), .Y(n4037) );
  AND2X1 U3696 ( .A(fifo_array[175]), .B(n5830), .Y(n363) );
  INVX1 U3697 ( .A(n363), .Y(n4038) );
  AND2X1 U3698 ( .A(fifo_array[147]), .B(n5832), .Y(n333) );
  INVX1 U3699 ( .A(n333), .Y(n4039) );
  AND2X1 U3700 ( .A(fifo_array[134]), .B(n5833), .Y(n320) );
  INVX1 U3701 ( .A(n320), .Y(n4040) );
  AND2X1 U3702 ( .A(fifo_array[126]), .B(n5833), .Y(n312) );
  INVX1 U3703 ( .A(n312), .Y(n4041) );
  AND2X1 U3704 ( .A(fifo_array[109]), .B(n5834), .Y(n293) );
  INVX1 U3705 ( .A(n293), .Y(n4042) );
  AND2X1 U3706 ( .A(fifo_array[97]), .B(n5835), .Y(n281) );
  INVX1 U3707 ( .A(n281), .Y(n4043) );
  AND2X1 U3708 ( .A(fifo_array[85]), .B(n5835), .Y(n269) );
  INVX1 U3709 ( .A(n269), .Y(n4044) );
  AND2X1 U3710 ( .A(fifo_array[68]), .B(n5836), .Y(n250) );
  INVX1 U3711 ( .A(n250), .Y(n4045) );
  AND2X1 U3712 ( .A(fifo_array[56]), .B(n5837), .Y(n238) );
  INVX1 U3713 ( .A(n238), .Y(n4046) );
  AND2X1 U3714 ( .A(fifo_array[44]), .B(n5836), .Y(n226) );
  INVX1 U3715 ( .A(n226), .Y(n4047) );
  AND2X1 U3716 ( .A(fifo_array[15]), .B(n5838), .Y(n194) );
  INVX1 U3717 ( .A(n194), .Y(n4048) );
  AND2X1 U3718 ( .A(fifo_array[3]), .B(n5839), .Y(n182) );
  INVX1 U3719 ( .A(n182), .Y(n4049) );
  INVX1 U3720 ( .A(n1635), .Y(n4050) );
  BUFX2 U3721 ( .A(n1634), .Y(n4051) );
  BUFX2 U3722 ( .A(n1637), .Y(n4052) );
  AND2X1 U3723 ( .A(n84), .B(n5773), .Y(n1584) );
  INVX1 U3724 ( .A(n1584), .Y(n4053) );
  AND2X1 U3725 ( .A(fifo_array[1331]), .B(n5776), .Y(n1553) );
  INVX1 U3726 ( .A(n1553), .Y(n4054) );
  AND2X1 U3727 ( .A(fifo_array[1322]), .B(n5777), .Y(n1544) );
  INVX1 U3728 ( .A(n1544), .Y(n4055) );
  AND2X1 U3729 ( .A(fifo_array[1309]), .B(n5777), .Y(n1531) );
  INVX1 U3730 ( .A(n1531), .Y(n4056) );
  AND2X1 U3731 ( .A(fifo_array[1288]), .B(n5778), .Y(n1509) );
  INVX1 U3732 ( .A(n1509), .Y(n4057) );
  AND2X1 U3733 ( .A(fifo_array[1279]), .B(n5779), .Y(n1500) );
  INVX1 U3734 ( .A(n1500), .Y(n4058) );
  AND2X1 U3735 ( .A(fifo_array[1266]), .B(n5779), .Y(n1487) );
  INVX1 U3736 ( .A(n1487), .Y(n4059) );
  AND2X1 U3737 ( .A(fifo_array[1243]), .B(n5781), .Y(n1463) );
  INVX1 U3738 ( .A(n1463), .Y(n4060) );
  AND2X1 U3739 ( .A(fifo_array[1231]), .B(n5780), .Y(n1451) );
  INVX1 U3740 ( .A(n1451), .Y(n4061) );
  AND2X1 U3741 ( .A(fifo_array[1219]), .B(n5781), .Y(n1439) );
  INVX1 U3742 ( .A(n1439), .Y(n4062) );
  AND2X1 U3743 ( .A(fifo_array[1197]), .B(n5783), .Y(n1416) );
  INVX1 U3744 ( .A(n1416), .Y(n4063) );
  AND2X1 U3745 ( .A(fifo_array[1184]), .B(n5782), .Y(n1403) );
  INVX1 U3746 ( .A(n1403), .Y(n4064) );
  AND2X1 U3747 ( .A(fifo_array[1176]), .B(n5783), .Y(n1395) );
  INVX1 U3748 ( .A(n1395), .Y(n4065) );
  AND2X1 U3749 ( .A(fifo_array[1149]), .B(n5784), .Y(n1367) );
  INVX1 U3750 ( .A(n1367), .Y(n4066) );
  AND2X1 U3751 ( .A(fifo_array[1137]), .B(n5785), .Y(n1355) );
  INVX1 U3752 ( .A(n1355), .Y(n4067) );
  AND2X1 U3753 ( .A(fifo_array[1118]), .B(n5786), .Y(n1335) );
  INVX1 U3754 ( .A(n1335), .Y(n4068) );
  AND2X1 U3755 ( .A(fifo_array[1106]), .B(n5786), .Y(n1323) );
  INVX1 U3756 ( .A(n1323), .Y(n4069) );
  AND2X1 U3757 ( .A(fifo_array[1094]), .B(n5787), .Y(n1311) );
  INVX1 U3758 ( .A(n1311), .Y(n4070) );
  AND2X1 U3759 ( .A(fifo_array[1083]), .B(n5788), .Y(n1299) );
  INVX1 U3760 ( .A(n1299), .Y(n4071) );
  AND2X1 U3761 ( .A(fifo_array[1044]), .B(n5791), .Y(n1258) );
  INVX1 U3762 ( .A(n1258), .Y(n4072) );
  AND2X1 U3763 ( .A(fifo_array[1030]), .B(n5790), .Y(n1244) );
  INVX1 U3764 ( .A(n1244), .Y(n4073) );
  AND2X1 U3765 ( .A(fifo_array[1018]), .B(n5791), .Y(n1232) );
  INVX1 U3766 ( .A(n1232), .Y(n4074) );
  AND2X1 U3767 ( .A(fifo_array[982]), .B(n5793), .Y(n1195) );
  INVX1 U3768 ( .A(n1195), .Y(n4075) );
  AND2X1 U3769 ( .A(fifo_array[975]), .B(n5793), .Y(n1188) );
  INVX1 U3770 ( .A(n1188), .Y(n4076) );
  AND2X1 U3771 ( .A(fifo_array[954]), .B(n5795), .Y(n1166) );
  INVX1 U3772 ( .A(n1166), .Y(n4077) );
  AND2X1 U3773 ( .A(fifo_array[948]), .B(n5794), .Y(n1160) );
  INVX1 U3774 ( .A(n1160), .Y(n4078) );
  AND2X1 U3775 ( .A(fifo_array[936]), .B(n5795), .Y(n1148) );
  INVX1 U3776 ( .A(n1148), .Y(n4079) );
  AND2X1 U3777 ( .A(fifo_array[921]), .B(n5796), .Y(n1132) );
  INVX1 U3778 ( .A(n1132), .Y(n4080) );
  AND2X1 U3779 ( .A(fifo_array[905]), .B(n5796), .Y(n1116) );
  INVX1 U3780 ( .A(n1116), .Y(n4081) );
  AND2X1 U3781 ( .A(fifo_array[893]), .B(n5797), .Y(n1104) );
  INVX1 U3782 ( .A(n1104), .Y(n4082) );
  AND2X1 U3783 ( .A(fifo_array[867]), .B(n5799), .Y(n1077) );
  INVX1 U3784 ( .A(n1077), .Y(n4083) );
  AND2X1 U3785 ( .A(fifo_array[858]), .B(n5798), .Y(n1068) );
  INVX1 U3786 ( .A(n1068), .Y(n4084) );
  AND2X1 U3787 ( .A(fifo_array[845]), .B(n5799), .Y(n1055) );
  INVX1 U3788 ( .A(n1055), .Y(n4085) );
  AND2X1 U3789 ( .A(fifo_array[815]), .B(n5801), .Y(n1024) );
  INVX1 U3790 ( .A(n1024), .Y(n4086) );
  AND2X1 U3791 ( .A(fifo_array[802]), .B(n5801), .Y(n1011) );
  INVX1 U3792 ( .A(n1011), .Y(n4087) );
  AND2X1 U3793 ( .A(fifo_array[785]), .B(n5803), .Y(n993) );
  INVX1 U3794 ( .A(n993), .Y(n4088) );
  AND2X1 U3795 ( .A(fifo_array[776]), .B(n5802), .Y(n984) );
  INVX1 U3796 ( .A(n984), .Y(n4089) );
  AND2X1 U3797 ( .A(fifo_array[763]), .B(n5802), .Y(n971) );
  INVX1 U3798 ( .A(n971), .Y(n4090) );
  AND2X1 U3799 ( .A(fifo_array[742]), .B(n5805), .Y(n949) );
  INVX1 U3800 ( .A(n949), .Y(n4091) );
  AND2X1 U3801 ( .A(fifo_array[733]), .B(n5804), .Y(n940) );
  INVX1 U3802 ( .A(n940), .Y(n4092) );
  AND2X1 U3803 ( .A(fifo_array[720]), .B(n5804), .Y(n927) );
  INVX1 U3804 ( .A(n927), .Y(n4093) );
  AND2X1 U3805 ( .A(fifo_array[697]), .B(n5806), .Y(n902) );
  INVX1 U3806 ( .A(n902), .Y(n4094) );
  AND2X1 U3807 ( .A(fifo_array[685]), .B(n5807), .Y(n890) );
  INVX1 U3808 ( .A(n890), .Y(n4095) );
  AND2X1 U3809 ( .A(fifo_array[673]), .B(n5807), .Y(n878) );
  INVX1 U3810 ( .A(n878), .Y(n4096) );
  AND2X1 U3811 ( .A(fifo_array[651]), .B(n5808), .Y(n855) );
  INVX1 U3812 ( .A(n855), .Y(n4097) );
  AND2X1 U3813 ( .A(fifo_array[638]), .B(n5809), .Y(n842) );
  INVX1 U3814 ( .A(n842), .Y(n4098) );
  AND2X1 U3815 ( .A(fifo_array[630]), .B(n5809), .Y(n834) );
  INVX1 U3816 ( .A(n834), .Y(n4099) );
  AND2X1 U3817 ( .A(fifo_array[603]), .B(n5811), .Y(n806) );
  INVX1 U3818 ( .A(n806), .Y(n4100) );
  AND2X1 U3819 ( .A(fifo_array[591]), .B(n5811), .Y(n794) );
  INVX1 U3820 ( .A(n794), .Y(n4101) );
  AND2X1 U3821 ( .A(fifo_array[572]), .B(n5812), .Y(n774) );
  INVX1 U3822 ( .A(n774), .Y(n4102) );
  AND2X1 U3823 ( .A(fifo_array[560]), .B(n5813), .Y(n762) );
  INVX1 U3824 ( .A(n762), .Y(n4103) );
  AND2X1 U3825 ( .A(fifo_array[548]), .B(n5813), .Y(n750) );
  INVX1 U3826 ( .A(n750), .Y(n4104) );
  AND2X1 U3827 ( .A(fifo_array[537]), .B(n5815), .Y(n738) );
  INVX1 U3828 ( .A(n738), .Y(n4105) );
  AND2X1 U3829 ( .A(fifo_array[498]), .B(n5817), .Y(n698) );
  INVX1 U3830 ( .A(n698), .Y(n4106) );
  AND2X1 U3831 ( .A(fifo_array[484]), .B(n5816), .Y(n684) );
  INVX1 U3832 ( .A(n684), .Y(n4107) );
  AND2X1 U3833 ( .A(fifo_array[472]), .B(n5817), .Y(n672) );
  INVX1 U3834 ( .A(n672), .Y(n4108) );
  AND2X1 U3835 ( .A(fifo_array[436]), .B(n5819), .Y(n635) );
  INVX1 U3836 ( .A(n635), .Y(n4109) );
  AND2X1 U3837 ( .A(fifo_array[429]), .B(n5819), .Y(n628) );
  INVX1 U3838 ( .A(n628), .Y(n4110) );
  AND2X1 U3839 ( .A(fifo_array[408]), .B(n5821), .Y(n606) );
  INVX1 U3840 ( .A(n606), .Y(n4111) );
  AND2X1 U3841 ( .A(fifo_array[402]), .B(n5820), .Y(n600) );
  INVX1 U3842 ( .A(n600), .Y(n4112) );
  AND2X1 U3843 ( .A(fifo_array[390]), .B(n5821), .Y(n588) );
  INVX1 U3844 ( .A(n588), .Y(n4113) );
  AND2X1 U3845 ( .A(fifo_array[375]), .B(n5822), .Y(n571) );
  INVX1 U3846 ( .A(n571), .Y(n4114) );
  AND2X1 U3847 ( .A(fifo_array[359]), .B(n5822), .Y(n555) );
  INVX1 U3848 ( .A(n555), .Y(n4115) );
  AND2X1 U3849 ( .A(fifo_array[347]), .B(n5823), .Y(n543) );
  INVX1 U3850 ( .A(n543), .Y(n4116) );
  AND2X1 U3851 ( .A(fifo_array[321]), .B(n5825), .Y(n515) );
  INVX1 U3852 ( .A(n515), .Y(n4117) );
  AND2X1 U3853 ( .A(fifo_array[312]), .B(n5824), .Y(n506) );
  INVX1 U3854 ( .A(n506), .Y(n4118) );
  AND2X1 U3855 ( .A(fifo_array[299]), .B(n5825), .Y(n493) );
  INVX1 U3856 ( .A(n493), .Y(n4119) );
  AND2X1 U3857 ( .A(fifo_array[269]), .B(n5827), .Y(n461) );
  INVX1 U3858 ( .A(n461), .Y(n4120) );
  AND2X1 U3859 ( .A(fifo_array[256]), .B(n5827), .Y(n448) );
  INVX1 U3860 ( .A(n448), .Y(n4121) );
  AND2X1 U3861 ( .A(fifo_array[239]), .B(n5829), .Y(n429) );
  INVX1 U3862 ( .A(n429), .Y(n4122) );
  AND2X1 U3863 ( .A(fifo_array[230]), .B(n5828), .Y(n420) );
  INVX1 U3864 ( .A(n420), .Y(n4123) );
  AND2X1 U3865 ( .A(fifo_array[217]), .B(n5828), .Y(n407) );
  INVX1 U3866 ( .A(n407), .Y(n4124) );
  AND2X1 U3867 ( .A(fifo_array[196]), .B(n5831), .Y(n384) );
  INVX1 U3868 ( .A(n384), .Y(n4125) );
  AND2X1 U3869 ( .A(fifo_array[187]), .B(n5830), .Y(n375) );
  INVX1 U3870 ( .A(n375), .Y(n4126) );
  AND2X1 U3871 ( .A(fifo_array[174]), .B(n5830), .Y(n362) );
  INVX1 U3872 ( .A(n362), .Y(n4127) );
  AND2X1 U3873 ( .A(fifo_array[151]), .B(n5832), .Y(n337) );
  INVX1 U3874 ( .A(n337), .Y(n4128) );
  AND2X1 U3875 ( .A(fifo_array[139]), .B(n5833), .Y(n325) );
  INVX1 U3876 ( .A(n325), .Y(n4129) );
  AND2X1 U3877 ( .A(fifo_array[127]), .B(n5833), .Y(n313) );
  INVX1 U3878 ( .A(n313), .Y(n4130) );
  AND2X1 U3879 ( .A(fifo_array[105]), .B(n5834), .Y(n289) );
  INVX1 U3880 ( .A(n289), .Y(n4131) );
  AND2X1 U3881 ( .A(fifo_array[92]), .B(n5835), .Y(n276) );
  INVX1 U3882 ( .A(n276), .Y(n4132) );
  AND2X1 U3883 ( .A(fifo_array[84]), .B(n5835), .Y(n268) );
  INVX1 U3884 ( .A(n268), .Y(n4133) );
  AND2X1 U3885 ( .A(fifo_array[57]), .B(n5837), .Y(n239) );
  INVX1 U3886 ( .A(n239), .Y(n4134) );
  AND2X1 U3887 ( .A(fifo_array[45]), .B(n5837), .Y(n227) );
  INVX1 U3888 ( .A(n227), .Y(n4135) );
  AND2X1 U3889 ( .A(fifo_array[26]), .B(n5838), .Y(n205) );
  INVX1 U3890 ( .A(n205), .Y(n4136) );
  AND2X1 U3891 ( .A(fifo_array[14]), .B(n5838), .Y(n193) );
  INVX1 U3892 ( .A(n193), .Y(n4137) );
  AND2X1 U3893 ( .A(fifo_array[2]), .B(n5839), .Y(n181) );
  INVX1 U3894 ( .A(n181), .Y(n4138) );
  OR2X1 U3895 ( .A(n103), .B(n5904), .Y(n1648) );
  INVX1 U3896 ( .A(n1648), .Y(n4139) );
  INVX1 U3897 ( .A(n1573), .Y(n4140) );
  AND2X1 U3898 ( .A(fifo_array[1319]), .B(n5776), .Y(n1541) );
  INVX1 U3899 ( .A(n1541), .Y(n4141) );
  AND2X1 U3900 ( .A(fifo_array[1306]), .B(n5777), .Y(n1528) );
  INVX1 U3901 ( .A(n1528), .Y(n4142) );
  AND2X1 U3902 ( .A(fifo_array[1287]), .B(n5778), .Y(n1508) );
  INVX1 U3903 ( .A(n1508), .Y(n4143) );
  AND2X1 U3904 ( .A(fifo_array[1278]), .B(n5778), .Y(n1499) );
  INVX1 U3905 ( .A(n1499), .Y(n4144) );
  AND2X1 U3906 ( .A(fifo_array[1265]), .B(n5779), .Y(n1486) );
  INVX1 U3907 ( .A(n1486), .Y(n4145) );
  AND2X1 U3908 ( .A(fifo_array[1244]), .B(n5780), .Y(n1464) );
  INVX1 U3909 ( .A(n1464), .Y(n4146) );
  AND2X1 U3910 ( .A(fifo_array[1232]), .B(n5780), .Y(n1452) );
  INVX1 U3911 ( .A(n1452), .Y(n4147) );
  AND2X1 U3912 ( .A(fifo_array[1220]), .B(n5781), .Y(n1440) );
  INVX1 U3913 ( .A(n1440), .Y(n4148) );
  AND2X1 U3914 ( .A(fifo_array[1191]), .B(n5782), .Y(n1410) );
  INVX1 U3915 ( .A(n1410), .Y(n4149) );
  AND2X1 U3916 ( .A(fifo_array[1179]), .B(n5783), .Y(n1398) );
  INVX1 U3917 ( .A(n1398), .Y(n4150) );
  AND2X1 U3918 ( .A(fifo_array[1155]), .B(n5785), .Y(n1373) );
  INVX1 U3919 ( .A(n1373), .Y(n4151) );
  AND2X1 U3920 ( .A(fifo_array[1142]), .B(n5784), .Y(n1360) );
  INVX1 U3921 ( .A(n1360), .Y(n4152) );
  AND2X1 U3922 ( .A(fifo_array[1134]), .B(n5785), .Y(n1352) );
  INVX1 U3923 ( .A(n1352), .Y(n4153) );
  AND2X1 U3924 ( .A(fifo_array[1117]), .B(n5787), .Y(n1334) );
  INVX1 U3925 ( .A(n1334), .Y(n4154) );
  AND2X1 U3926 ( .A(fifo_array[1105]), .B(n5786), .Y(n1322) );
  INVX1 U3927 ( .A(n1322), .Y(n4155) );
  AND2X1 U3928 ( .A(fifo_array[1093]), .B(n5787), .Y(n1310) );
  INVX1 U3929 ( .A(n1310), .Y(n4156) );
  AND2X1 U3930 ( .A(fifo_array[1088]), .B(n5789), .Y(n1304) );
  INVX1 U3931 ( .A(n1304), .Y(n4157) );
  AND2X1 U3932 ( .A(fifo_array[1082]), .B(n5789), .Y(n1298) );
  INVX1 U3933 ( .A(n1298), .Y(n4158) );
  AND2X1 U3934 ( .A(fifo_array[1047]), .B(n5791), .Y(n1261) );
  INVX1 U3935 ( .A(n1261), .Y(n4159) );
  AND2X1 U3936 ( .A(fifo_array[1031]), .B(n5790), .Y(n1245) );
  INVX1 U3937 ( .A(n1245), .Y(n4160) );
  AND2X1 U3938 ( .A(fifo_array[1019]), .B(n5790), .Y(n1233) );
  INVX1 U3939 ( .A(n1233), .Y(n4161) );
  AND2X1 U3940 ( .A(fifo_array[996]), .B(n5793), .Y(n1209) );
  INVX1 U3941 ( .A(n1209), .Y(n4162) );
  AND2X1 U3942 ( .A(fifo_array[990]), .B(n5792), .Y(n1203) );
  INVX1 U3943 ( .A(n1203), .Y(n4163) );
  AND2X1 U3944 ( .A(fifo_array[978]), .B(n5793), .Y(n1191) );
  INVX1 U3945 ( .A(n1191), .Y(n4164) );
  AND2X1 U3946 ( .A(fifo_array[940]), .B(n5795), .Y(n1152) );
  INVX1 U3947 ( .A(n1152), .Y(n4165) );
  AND2X1 U3948 ( .A(fifo_array[933]), .B(n5795), .Y(n1145) );
  INVX1 U3949 ( .A(n1145), .Y(n4166) );
  AND2X1 U3950 ( .A(fifo_array[918]), .B(n5797), .Y(n1129) );
  INVX1 U3951 ( .A(n1129), .Y(n4167) );
  AND2X1 U3952 ( .A(fifo_array[904]), .B(n5796), .Y(n1115) );
  INVX1 U3953 ( .A(n1115), .Y(n4168) );
  AND2X1 U3954 ( .A(fifo_array[892]), .B(n5797), .Y(n1103) );
  INVX1 U3955 ( .A(n1103), .Y(n4169) );
  AND2X1 U3956 ( .A(fifo_array[868]), .B(n5799), .Y(n1078) );
  INVX1 U3957 ( .A(n1078), .Y(n4170) );
  AND2X1 U3958 ( .A(fifo_array[859]), .B(n5798), .Y(n1069) );
  INVX1 U3959 ( .A(n1069), .Y(n4171) );
  AND2X1 U3960 ( .A(fifo_array[846]), .B(n5798), .Y(n1056) );
  INVX1 U3961 ( .A(n1056), .Y(n4172) );
  AND2X1 U3962 ( .A(fifo_array[827]), .B(n5801), .Y(n1036) );
  INVX1 U3963 ( .A(n1036), .Y(n4173) );
  AND2X1 U3964 ( .A(fifo_array[818]), .B(n5800), .Y(n1027) );
  INVX1 U3965 ( .A(n1027), .Y(n4174) );
  AND2X1 U3966 ( .A(fifo_array[805]), .B(n5800), .Y(n1014) );
  INVX1 U3967 ( .A(n1014), .Y(n4175) );
  AND2X1 U3968 ( .A(fifo_array[773]), .B(n5803), .Y(n981) );
  INVX1 U3969 ( .A(n981), .Y(n4176) );
  AND2X1 U3970 ( .A(fifo_array[760]), .B(n5802), .Y(n968) );
  INVX1 U3971 ( .A(n968), .Y(n4177) );
  AND2X1 U3972 ( .A(fifo_array[741]), .B(n5805), .Y(n948) );
  INVX1 U3973 ( .A(n948), .Y(n4178) );
  AND2X1 U3974 ( .A(fifo_array[732]), .B(n5804), .Y(n939) );
  INVX1 U3975 ( .A(n939), .Y(n4179) );
  AND2X1 U3976 ( .A(fifo_array[719]), .B(n5804), .Y(n926) );
  INVX1 U3977 ( .A(n926), .Y(n4180) );
  AND2X1 U3978 ( .A(fifo_array[698]), .B(n5806), .Y(n903) );
  INVX1 U3979 ( .A(n903), .Y(n4181) );
  AND2X1 U3980 ( .A(fifo_array[686]), .B(n5807), .Y(n891) );
  INVX1 U3981 ( .A(n891), .Y(n4182) );
  AND2X1 U3982 ( .A(fifo_array[674]), .B(n5806), .Y(n879) );
  INVX1 U3983 ( .A(n879), .Y(n4183) );
  AND2X1 U3984 ( .A(fifo_array[645]), .B(n5809), .Y(n849) );
  INVX1 U3985 ( .A(n849), .Y(n4184) );
  AND2X1 U3986 ( .A(fifo_array[633]), .B(n5808), .Y(n837) );
  INVX1 U3987 ( .A(n837), .Y(n4185) );
  AND2X1 U3988 ( .A(fifo_array[609]), .B(n5810), .Y(n812) );
  INVX1 U3989 ( .A(n812), .Y(n4186) );
  AND2X1 U3990 ( .A(fifo_array[596]), .B(n5811), .Y(n799) );
  INVX1 U3991 ( .A(n799), .Y(n4187) );
  AND2X1 U3992 ( .A(fifo_array[588]), .B(n5811), .Y(n791) );
  INVX1 U3993 ( .A(n791), .Y(n4188) );
  AND2X1 U3994 ( .A(fifo_array[571]), .B(n5812), .Y(n773) );
  INVX1 U3995 ( .A(n773), .Y(n4189) );
  AND2X1 U3996 ( .A(fifo_array[559]), .B(n5813), .Y(n761) );
  INVX1 U3997 ( .A(n761), .Y(n4190) );
  AND2X1 U3998 ( .A(fifo_array[547]), .B(n5813), .Y(n749) );
  INVX1 U3999 ( .A(n749), .Y(n4191) );
  AND2X1 U4000 ( .A(fifo_array[542]), .B(n5815), .Y(n743) );
  INVX1 U4001 ( .A(n743), .Y(n4192) );
  AND2X1 U4002 ( .A(fifo_array[536]), .B(n5815), .Y(n737) );
  INVX1 U4003 ( .A(n737), .Y(n4193) );
  AND2X1 U4004 ( .A(fifo_array[501]), .B(n5816), .Y(n701) );
  INVX1 U4005 ( .A(n701), .Y(n4194) );
  AND2X1 U4006 ( .A(fifo_array[485]), .B(n5816), .Y(n685) );
  INVX1 U4007 ( .A(n685), .Y(n4195) );
  AND2X1 U4008 ( .A(fifo_array[473]), .B(n5817), .Y(n673) );
  INVX1 U4009 ( .A(n673), .Y(n4196) );
  AND2X1 U4010 ( .A(fifo_array[450]), .B(n5819), .Y(n649) );
  INVX1 U4011 ( .A(n649), .Y(n4197) );
  AND2X1 U4012 ( .A(fifo_array[444]), .B(n5818), .Y(n643) );
  INVX1 U4013 ( .A(n643), .Y(n4198) );
  AND2X1 U4014 ( .A(fifo_array[432]), .B(n5819), .Y(n631) );
  INVX1 U4015 ( .A(n631), .Y(n4199) );
  AND2X1 U4016 ( .A(fifo_array[394]), .B(n5821), .Y(n592) );
  INVX1 U4017 ( .A(n592), .Y(n4200) );
  AND2X1 U4018 ( .A(fifo_array[387]), .B(n5821), .Y(n585) );
  INVX1 U4019 ( .A(n585), .Y(n4201) );
  AND2X1 U4020 ( .A(fifo_array[372]), .B(n5823), .Y(n568) );
  INVX1 U4021 ( .A(n568), .Y(n4202) );
  AND2X1 U4022 ( .A(fifo_array[358]), .B(n5822), .Y(n554) );
  INVX1 U4023 ( .A(n554), .Y(n4203) );
  AND2X1 U4024 ( .A(fifo_array[346]), .B(n5823), .Y(n542) );
  INVX1 U4025 ( .A(n542), .Y(n4204) );
  AND2X1 U4026 ( .A(fifo_array[322]), .B(n5825), .Y(n516) );
  INVX1 U4027 ( .A(n516), .Y(n4205) );
  AND2X1 U4028 ( .A(fifo_array[313]), .B(n5824), .Y(n507) );
  INVX1 U4029 ( .A(n507), .Y(n4206) );
  AND2X1 U4030 ( .A(fifo_array[300]), .B(n5824), .Y(n494) );
  INVX1 U4031 ( .A(n494), .Y(n4207) );
  AND2X1 U4032 ( .A(fifo_array[281]), .B(n5827), .Y(n473) );
  INVX1 U4033 ( .A(n473), .Y(n4208) );
  AND2X1 U4034 ( .A(fifo_array[272]), .B(n5826), .Y(n464) );
  INVX1 U4035 ( .A(n464), .Y(n4209) );
  AND2X1 U4036 ( .A(fifo_array[259]), .B(n5826), .Y(n451) );
  INVX1 U4037 ( .A(n451), .Y(n4210) );
  AND2X1 U4038 ( .A(fifo_array[227]), .B(n5829), .Y(n417) );
  INVX1 U4039 ( .A(n417), .Y(n4211) );
  AND2X1 U4040 ( .A(fifo_array[214]), .B(n5828), .Y(n404) );
  INVX1 U4041 ( .A(n404), .Y(n4212) );
  AND2X1 U4042 ( .A(fifo_array[195]), .B(n5831), .Y(n383) );
  INVX1 U4043 ( .A(n383), .Y(n4213) );
  AND2X1 U4044 ( .A(fifo_array[186]), .B(n5830), .Y(n374) );
  INVX1 U4045 ( .A(n374), .Y(n4214) );
  AND2X1 U4046 ( .A(fifo_array[173]), .B(n5830), .Y(n361) );
  INVX1 U4047 ( .A(n361), .Y(n4215) );
  AND2X1 U4048 ( .A(fifo_array[152]), .B(n5832), .Y(n338) );
  INVX1 U4049 ( .A(n338), .Y(n4216) );
  AND2X1 U4050 ( .A(fifo_array[140]), .B(n5833), .Y(n326) );
  INVX1 U4051 ( .A(n326), .Y(n4217) );
  AND2X1 U4052 ( .A(fifo_array[128]), .B(n5832), .Y(n314) );
  INVX1 U4053 ( .A(n314), .Y(n4218) );
  AND2X1 U4054 ( .A(fifo_array[99]), .B(n5835), .Y(n283) );
  INVX1 U4055 ( .A(n283), .Y(n4219) );
  AND2X1 U4056 ( .A(fifo_array[87]), .B(n5834), .Y(n271) );
  INVX1 U4057 ( .A(n271), .Y(n4220) );
  AND2X1 U4058 ( .A(fifo_array[63]), .B(n5836), .Y(n245) );
  INVX1 U4059 ( .A(n245), .Y(n4221) );
  AND2X1 U4060 ( .A(fifo_array[50]), .B(n5837), .Y(n232) );
  INVX1 U4061 ( .A(n232), .Y(n4222) );
  AND2X1 U4062 ( .A(fifo_array[42]), .B(n5837), .Y(n224) );
  INVX1 U4063 ( .A(n224), .Y(n4223) );
  AND2X1 U4064 ( .A(fifo_array[25]), .B(n5838), .Y(n204) );
  INVX1 U4065 ( .A(n204), .Y(n4224) );
  AND2X1 U4066 ( .A(fifo_array[13]), .B(n5839), .Y(n192) );
  INVX1 U4067 ( .A(n192), .Y(n4225) );
  AND2X1 U4068 ( .A(fifo_array[1]), .B(n5839), .Y(n180) );
  INVX1 U4069 ( .A(n180), .Y(n4226) );
  AND2X1 U4070 ( .A(fillcount[2]), .B(fillcount[3]), .Y(n1650) );
  INVX1 U4071 ( .A(n1650), .Y(n4227) );
  AND2X1 U4072 ( .A(put), .B(n5895), .Y(n1647) );
  INVX1 U4073 ( .A(n1647), .Y(n4228) );
  AND2X1 U4074 ( .A(n5846), .B(n5851), .Y(n5847) );
  INVX1 U4075 ( .A(n5847), .Y(n4229) );
  AND2X1 U4076 ( .A(n4323), .B(n5845), .Y(n1583) );
  INVX1 U4077 ( .A(n1583), .Y(n4230) );
  INVX1 U4078 ( .A(n1568), .Y(n4231) );
  AND2X1 U4079 ( .A(fifo_array[1329]), .B(n5776), .Y(n1551) );
  INVX1 U4080 ( .A(n1551), .Y(n4232) );
  AND2X1 U4081 ( .A(fifo_array[1320]), .B(n5776), .Y(n1542) );
  INVX1 U4082 ( .A(n1542), .Y(n4233) );
  AND2X1 U4083 ( .A(fifo_array[1307]), .B(n5777), .Y(n1529) );
  INVX1 U4084 ( .A(n1529), .Y(n4234) );
  AND2X1 U4085 ( .A(fifo_array[1277]), .B(n5778), .Y(n1498) );
  INVX1 U4086 ( .A(n1498), .Y(n4235) );
  AND2X1 U4087 ( .A(fifo_array[1264]), .B(n5779), .Y(n1485) );
  INVX1 U4088 ( .A(n1485), .Y(n4236) );
  AND2X1 U4089 ( .A(fifo_array[1233]), .B(n5780), .Y(n1453) );
  INVX1 U4090 ( .A(n1453), .Y(n4237) );
  AND2X1 U4091 ( .A(fifo_array[1221]), .B(n5781), .Y(n1441) );
  INVX1 U4092 ( .A(n1441), .Y(n4238) );
  AND2X1 U4093 ( .A(fifo_array[1202]), .B(n5782), .Y(n1421) );
  INVX1 U4094 ( .A(n1421), .Y(n4239) );
  AND2X1 U4095 ( .A(fifo_array[1190]), .B(n5782), .Y(n1409) );
  INVX1 U4096 ( .A(n1409), .Y(n4240) );
  AND2X1 U4097 ( .A(fifo_array[1178]), .B(n5783), .Y(n1397) );
  INVX1 U4098 ( .A(n1397), .Y(n4241) );
  AND2X1 U4099 ( .A(fifo_array[1159]), .B(n5784), .Y(n1377) );
  INVX1 U4100 ( .A(n1377), .Y(n4242) );
  AND2X1 U4101 ( .A(fifo_array[1147]), .B(n5784), .Y(n1365) );
  INVX1 U4102 ( .A(n1365), .Y(n4243) );
  AND2X1 U4103 ( .A(fifo_array[1135]), .B(n5785), .Y(n1353) );
  INVX1 U4104 ( .A(n1353), .Y(n4244) );
  AND2X1 U4105 ( .A(fifo_array[1113]), .B(n5786), .Y(n1330) );
  INVX1 U4106 ( .A(n1330), .Y(n4245) );
  AND2X1 U4107 ( .A(fifo_array[1100]), .B(n5786), .Y(n1317) );
  INVX1 U4108 ( .A(n1317), .Y(n4246) );
  AND2X1 U4109 ( .A(fifo_array[1092]), .B(n5787), .Y(n1309) );
  INVX1 U4110 ( .A(n1309), .Y(n4247) );
  AND2X1 U4111 ( .A(fifo_array[1087]), .B(n5789), .Y(n1303) );
  INVX1 U4112 ( .A(n1303), .Y(n4248) );
  AND2X1 U4113 ( .A(fifo_array[1081]), .B(n5788), .Y(n1297) );
  INVX1 U4114 ( .A(n1297), .Y(n4249) );
  AND2X1 U4115 ( .A(fifo_array[1038]), .B(n5790), .Y(n1252) );
  INVX1 U4116 ( .A(n1252), .Y(n4250) );
  AND2X1 U4117 ( .A(fifo_array[1032]), .B(n5791), .Y(n1246) );
  INVX1 U4118 ( .A(n1246), .Y(n4251) );
  AND2X1 U4119 ( .A(fifo_array[1020]), .B(n5791), .Y(n1234) );
  INVX1 U4120 ( .A(n1234), .Y(n4252) );
  AND2X1 U4121 ( .A(fifo_array[1005]), .B(n5792), .Y(n1218) );
  INVX1 U4122 ( .A(n1218), .Y(n4253) );
  AND2X1 U4123 ( .A(fifo_array[989]), .B(n5792), .Y(n1202) );
  INVX1 U4124 ( .A(n1202), .Y(n4254) );
  AND2X1 U4125 ( .A(fifo_array[977]), .B(n5793), .Y(n1190) );
  INVX1 U4126 ( .A(n1190), .Y(n4255) );
  AND2X1 U4127 ( .A(fifo_array[960]), .B(n5794), .Y(n1172) );
  INVX1 U4128 ( .A(n1172), .Y(n4256) );
  AND2X1 U4129 ( .A(fifo_array[946]), .B(n5794), .Y(n1158) );
  INVX1 U4130 ( .A(n1158), .Y(n4257) );
  AND2X1 U4131 ( .A(fifo_array[934]), .B(n5795), .Y(n1146) );
  INVX1 U4132 ( .A(n1146), .Y(n4258) );
  AND2X1 U4133 ( .A(fifo_array[898]), .B(n5796), .Y(n1109) );
  INVX1 U4134 ( .A(n1109), .Y(n4259) );
  AND2X1 U4135 ( .A(fifo_array[891]), .B(n5797), .Y(n1102) );
  INVX1 U4136 ( .A(n1102), .Y(n4260) );
  AND2X1 U4137 ( .A(fifo_array[869]), .B(n5799), .Y(n1079) );
  INVX1 U4138 ( .A(n1079), .Y(n4261) );
  AND2X1 U4139 ( .A(fifo_array[860]), .B(n5798), .Y(n1070) );
  INVX1 U4140 ( .A(n1070), .Y(n4262) );
  AND2X1 U4141 ( .A(fifo_array[847]), .B(n5798), .Y(n1057) );
  INVX1 U4142 ( .A(n1057), .Y(n4263) );
  AND2X1 U4143 ( .A(fifo_array[826]), .B(n5801), .Y(n1035) );
  INVX1 U4144 ( .A(n1035), .Y(n4264) );
  AND2X1 U4145 ( .A(fifo_array[817]), .B(n5800), .Y(n1026) );
  INVX1 U4146 ( .A(n1026), .Y(n4265) );
  AND2X1 U4147 ( .A(fifo_array[804]), .B(n5800), .Y(n1013) );
  INVX1 U4148 ( .A(n1013), .Y(n4266) );
  AND2X1 U4149 ( .A(fifo_array[783]), .B(n5803), .Y(n991) );
  INVX1 U4150 ( .A(n991), .Y(n4267) );
  AND2X1 U4151 ( .A(fifo_array[774]), .B(n5802), .Y(n982) );
  INVX1 U4152 ( .A(n982), .Y(n4268) );
  AND2X1 U4153 ( .A(fifo_array[761]), .B(n5803), .Y(n969) );
  INVX1 U4154 ( .A(n969), .Y(n4269) );
  AND2X1 U4155 ( .A(fifo_array[731]), .B(n5805), .Y(n938) );
  INVX1 U4156 ( .A(n938), .Y(n4270) );
  AND2X1 U4157 ( .A(fifo_array[718]), .B(n5805), .Y(n925) );
  INVX1 U4158 ( .A(n925), .Y(n4271) );
  AND2X1 U4159 ( .A(fifo_array[687]), .B(n5807), .Y(n892) );
  INVX1 U4160 ( .A(n892), .Y(n4272) );
  AND2X1 U4161 ( .A(fifo_array[675]), .B(n5807), .Y(n880) );
  INVX1 U4162 ( .A(n880), .Y(n4273) );
  AND2X1 U4163 ( .A(fifo_array[656]), .B(n5808), .Y(n860) );
  INVX1 U4164 ( .A(n860), .Y(n4274) );
  AND2X1 U4165 ( .A(fifo_array[644]), .B(n5809), .Y(n848) );
  INVX1 U4166 ( .A(n848), .Y(n4275) );
  AND2X1 U4167 ( .A(fifo_array[632]), .B(n5809), .Y(n836) );
  INVX1 U4168 ( .A(n836), .Y(n4276) );
  AND2X1 U4169 ( .A(fifo_array[613]), .B(n5810), .Y(n816) );
  INVX1 U4170 ( .A(n816), .Y(n4277) );
  AND2X1 U4171 ( .A(fifo_array[601]), .B(n5811), .Y(n804) );
  INVX1 U4172 ( .A(n804), .Y(n4278) );
  AND2X1 U4173 ( .A(fifo_array[589]), .B(n5811), .Y(n792) );
  INVX1 U4174 ( .A(n792), .Y(n4279) );
  AND2X1 U4175 ( .A(fifo_array[567]), .B(n5812), .Y(n769) );
  INVX1 U4176 ( .A(n769), .Y(n4280) );
  AND2X1 U4177 ( .A(fifo_array[554]), .B(n5813), .Y(n756) );
  INVX1 U4178 ( .A(n756), .Y(n4281) );
  AND2X1 U4179 ( .A(fifo_array[546]), .B(n5813), .Y(n748) );
  INVX1 U4180 ( .A(n748), .Y(n4282) );
  AND2X1 U4181 ( .A(fifo_array[541]), .B(n5814), .Y(n742) );
  INVX1 U4182 ( .A(n742), .Y(n4283) );
  AND2X1 U4183 ( .A(fifo_array[535]), .B(n5815), .Y(n736) );
  INVX1 U4184 ( .A(n736), .Y(n4284) );
  AND2X1 U4185 ( .A(fifo_array[492]), .B(n5817), .Y(n692) );
  INVX1 U4186 ( .A(n692), .Y(n4285) );
  AND2X1 U4187 ( .A(fifo_array[486]), .B(n5816), .Y(n686) );
  INVX1 U4188 ( .A(n686), .Y(n4286) );
  AND2X1 U4189 ( .A(fifo_array[474]), .B(n5817), .Y(n674) );
  INVX1 U4190 ( .A(n674), .Y(n4287) );
  AND2X1 U4191 ( .A(fifo_array[459]), .B(n5818), .Y(n658) );
  INVX1 U4192 ( .A(n658), .Y(n4288) );
  AND2X1 U4193 ( .A(fifo_array[443]), .B(n5818), .Y(n642) );
  INVX1 U4194 ( .A(n642), .Y(n4289) );
  AND2X1 U4195 ( .A(fifo_array[431]), .B(n5819), .Y(n630) );
  INVX1 U4196 ( .A(n630), .Y(n4290) );
  AND2X1 U4197 ( .A(fifo_array[414]), .B(n5820), .Y(n612) );
  INVX1 U4198 ( .A(n612), .Y(n4291) );
  AND2X1 U4199 ( .A(fifo_array[400]), .B(n5820), .Y(n598) );
  INVX1 U4200 ( .A(n598), .Y(n4292) );
  AND2X1 U4201 ( .A(fifo_array[388]), .B(n5821), .Y(n586) );
  INVX1 U4202 ( .A(n586), .Y(n4293) );
  AND2X1 U4203 ( .A(fifo_array[352]), .B(n5822), .Y(n548) );
  INVX1 U4204 ( .A(n548), .Y(n4294) );
  AND2X1 U4205 ( .A(fifo_array[345]), .B(n5823), .Y(n541) );
  INVX1 U4206 ( .A(n541), .Y(n4295) );
  AND2X1 U4207 ( .A(fifo_array[323]), .B(n5825), .Y(n517) );
  INVX1 U4208 ( .A(n517), .Y(n4296) );
  AND2X1 U4209 ( .A(fifo_array[314]), .B(n5824), .Y(n508) );
  INVX1 U4210 ( .A(n508), .Y(n4297) );
  AND2X1 U4211 ( .A(fifo_array[301]), .B(n5824), .Y(n495) );
  INVX1 U4212 ( .A(n495), .Y(n4298) );
  AND2X1 U4213 ( .A(fifo_array[280]), .B(n5827), .Y(n472) );
  INVX1 U4214 ( .A(n472), .Y(n4299) );
  AND2X1 U4215 ( .A(fifo_array[271]), .B(n5826), .Y(n463) );
  INVX1 U4216 ( .A(n463), .Y(n4300) );
  AND2X1 U4217 ( .A(fifo_array[258]), .B(n5826), .Y(n450) );
  INVX1 U4218 ( .A(n450), .Y(n4301) );
  AND2X1 U4219 ( .A(fifo_array[237]), .B(n5829), .Y(n427) );
  INVX1 U4220 ( .A(n427), .Y(n4302) );
  AND2X1 U4221 ( .A(fifo_array[228]), .B(n5828), .Y(n418) );
  INVX1 U4222 ( .A(n418), .Y(n4303) );
  AND2X1 U4223 ( .A(fifo_array[215]), .B(n5829), .Y(n405) );
  INVX1 U4224 ( .A(n405), .Y(n4304) );
  AND2X1 U4225 ( .A(fifo_array[185]), .B(n5831), .Y(n373) );
  INVX1 U4226 ( .A(n373), .Y(n4305) );
  AND2X1 U4227 ( .A(fifo_array[172]), .B(n5831), .Y(n360) );
  INVX1 U4228 ( .A(n360), .Y(n4306) );
  AND2X1 U4229 ( .A(fifo_array[141]), .B(n5833), .Y(n327) );
  INVX1 U4230 ( .A(n327), .Y(n4307) );
  AND2X1 U4231 ( .A(fifo_array[129]), .B(n5833), .Y(n315) );
  INVX1 U4232 ( .A(n315), .Y(n4308) );
  AND2X1 U4233 ( .A(fifo_array[110]), .B(n5834), .Y(n294) );
  INVX1 U4234 ( .A(n294), .Y(n4309) );
  AND2X1 U4235 ( .A(fifo_array[98]), .B(n5835), .Y(n282) );
  INVX1 U4236 ( .A(n282), .Y(n4310) );
  AND2X1 U4237 ( .A(fifo_array[86]), .B(n5835), .Y(n270) );
  INVX1 U4238 ( .A(n270), .Y(n4311) );
  AND2X1 U4239 ( .A(fifo_array[67]), .B(n5836), .Y(n249) );
  INVX1 U4240 ( .A(n249), .Y(n4312) );
  AND2X1 U4241 ( .A(fifo_array[55]), .B(n5837), .Y(n237) );
  INVX1 U4242 ( .A(n237), .Y(n4313) );
  AND2X1 U4243 ( .A(fifo_array[43]), .B(n5837), .Y(n225) );
  INVX1 U4244 ( .A(n225), .Y(n4314) );
  AND2X1 U4245 ( .A(fifo_array[21]), .B(n5838), .Y(n200) );
  INVX1 U4246 ( .A(n200), .Y(n4315) );
  AND2X1 U4247 ( .A(fifo_array[8]), .B(n5838), .Y(n187) );
  INVX1 U4248 ( .A(n187), .Y(n4316) );
  AND2X1 U4249 ( .A(fifo_array[0]), .B(n5839), .Y(n179) );
  INVX1 U4250 ( .A(n179), .Y(n4317) );
  AND2X1 U4251 ( .A(n5903), .B(n5896), .Y(n1640) );
  INVX1 U4252 ( .A(n1640), .Y(n4318) );
  AND2X1 U4253 ( .A(n5904), .B(n103), .Y(n5846) );
  INVX1 U4254 ( .A(n5846), .Y(n4319) );
  AND2X1 U4255 ( .A(n5847), .B(n5850), .Y(n5848) );
  INVX1 U4256 ( .A(n5848), .Y(n4320) );
  BUFX2 U4257 ( .A(n1632), .Y(n4321) );
  AND2X1 U4258 ( .A(n1568), .B(n5845), .Y(n1566) );
  INVX1 U4259 ( .A(n1566), .Y(n4322) );
  INVX1 U4260 ( .A(n5634), .Y(n5691) );
  INVX1 U4261 ( .A(n5634), .Y(n5690) );
  INVX1 U4262 ( .A(n5633), .Y(n5689) );
  INVX1 U4263 ( .A(n5626), .Y(n5688) );
  INVX1 U4264 ( .A(n5631), .Y(n5687) );
  INVX1 U4265 ( .A(n5626), .Y(n5686) );
  INVX1 U4266 ( .A(n5626), .Y(n5685) );
  INVX1 U4267 ( .A(n5626), .Y(n5684) );
  INVX1 U4268 ( .A(n5626), .Y(n5683) );
  INVX1 U4269 ( .A(n5626), .Y(n5682) );
  INVX1 U4270 ( .A(n5632), .Y(n5681) );
  INVX1 U4271 ( .A(n5633), .Y(n5680) );
  INVX1 U4272 ( .A(n5627), .Y(n5679) );
  INVX1 U4273 ( .A(n5627), .Y(n5678) );
  INVX1 U4274 ( .A(n5627), .Y(n5677) );
  INVX1 U4275 ( .A(n5629), .Y(n5676) );
  INVX1 U4276 ( .A(n5630), .Y(n5675) );
  INVX1 U4277 ( .A(n5628), .Y(n5674) );
  INVX1 U4278 ( .A(n5628), .Y(n5673) );
  INVX1 U4279 ( .A(n5628), .Y(n5672) );
  INVX1 U4280 ( .A(n5628), .Y(n5671) );
  INVX1 U4281 ( .A(n5629), .Y(n5670) );
  INVX1 U4282 ( .A(n5629), .Y(n5669) );
  INVX1 U4283 ( .A(n5629), .Y(n5668) );
  INVX1 U4284 ( .A(n5630), .Y(n5667) );
  INVX1 U4285 ( .A(n5630), .Y(n5666) );
  INVX1 U4286 ( .A(n5630), .Y(n5665) );
  INVX1 U4287 ( .A(n5632), .Y(n5664) );
  INVX1 U4288 ( .A(n5634), .Y(n5663) );
  INVX1 U4289 ( .A(n5633), .Y(n5662) );
  INVX1 U4290 ( .A(n5631), .Y(n5661) );
  INVX1 U4291 ( .A(n5631), .Y(n5660) );
  INVX1 U4292 ( .A(n5632), .Y(n5659) );
  INVX1 U4293 ( .A(n5631), .Y(n5658) );
  INVX1 U4294 ( .A(n5631), .Y(n5657) );
  INVX1 U4295 ( .A(n5631), .Y(n5656) );
  INVX1 U4296 ( .A(n5632), .Y(n5655) );
  INVX1 U4297 ( .A(n5632), .Y(n5654) );
  INVX1 U4298 ( .A(n5632), .Y(n5653) );
  INVX1 U4299 ( .A(n5633), .Y(n5652) );
  INVX1 U4300 ( .A(n5633), .Y(n5651) );
  INVX1 U4301 ( .A(n5633), .Y(n5650) );
  INVX1 U4302 ( .A(n5634), .Y(n5649) );
  INVX1 U4303 ( .A(n5634), .Y(n5648) );
  INVX1 U4304 ( .A(n5634), .Y(n5647) );
  INVX1 U4305 ( .A(n5635), .Y(n5646) );
  INVX1 U4306 ( .A(n5635), .Y(n5645) );
  INVX1 U4307 ( .A(n5635), .Y(n5644) );
  INVX1 U4308 ( .A(n5636), .Y(n5643) );
  INVX1 U4309 ( .A(n5636), .Y(n5642) );
  INVX1 U4310 ( .A(n5636), .Y(n5641) );
  INVX1 U4311 ( .A(n5637), .Y(n5640) );
  INVX1 U4312 ( .A(n5637), .Y(n5639) );
  INVX1 U4313 ( .A(n5637), .Y(n5638) );
  INVX1 U4314 ( .A(n5636), .Y(n5693) );
  INVX1 U4315 ( .A(n5637), .Y(n5692) );
  INVX1 U4316 ( .A(n5695), .Y(n5626) );
  INVX1 U4317 ( .A(n5695), .Y(n5627) );
  INVX1 U4318 ( .A(n5694), .Y(n5628) );
  INVX1 U4319 ( .A(n5694), .Y(n5629) );
  INVX1 U4320 ( .A(n5694), .Y(n5630) );
  INVX1 U4321 ( .A(n5695), .Y(n5631) );
  INVX1 U4322 ( .A(n5695), .Y(n5632) );
  INVX1 U4323 ( .A(n5695), .Y(n5633) );
  INVX1 U4324 ( .A(n5695), .Y(n5634) );
  INVX1 U4325 ( .A(n5843), .Y(n5722) );
  INVX1 U4326 ( .A(n5843), .Y(n5721) );
  INVX1 U4327 ( .A(n5843), .Y(n5720) );
  INVX1 U4328 ( .A(n5843), .Y(n5719) );
  INVX1 U4329 ( .A(n5843), .Y(n5718) );
  INVX1 U4330 ( .A(n5843), .Y(n5717) );
  INVX1 U4331 ( .A(n5843), .Y(n5716) );
  INVX1 U4332 ( .A(n5843), .Y(n5715) );
  INVX1 U4333 ( .A(n5843), .Y(n5714) );
  INVX1 U4334 ( .A(n5843), .Y(n5713) );
  INVX1 U4335 ( .A(n5843), .Y(n5712) );
  INVX1 U4336 ( .A(n5843), .Y(n5711) );
  INVX1 U4337 ( .A(n5843), .Y(n5710) );
  INVX1 U4338 ( .A(n5843), .Y(n5709) );
  INVX1 U4339 ( .A(n5843), .Y(n5708) );
  INVX1 U4340 ( .A(n5843), .Y(n5707) );
  INVX1 U4341 ( .A(n5843), .Y(n5706) );
  INVX1 U4342 ( .A(n5843), .Y(n5705) );
  INVX1 U4343 ( .A(n5842), .Y(n5729) );
  INVX1 U4344 ( .A(n5842), .Y(n5728) );
  INVX1 U4345 ( .A(n5842), .Y(n5727) );
  INVX1 U4346 ( .A(n5842), .Y(n5726) );
  INVX1 U4347 ( .A(n5842), .Y(n5725) );
  INVX1 U4348 ( .A(n5842), .Y(n5724) );
  INVX1 U4349 ( .A(n5842), .Y(n5730) );
  INVX1 U4350 ( .A(n4323), .Y(n5773) );
  INVX1 U4351 ( .A(n1523), .Y(n5776) );
  INVX1 U4352 ( .A(n1523), .Y(n5777) );
  INVX1 U4353 ( .A(n5844), .Y(n5694) );
  INVX1 U4354 ( .A(n5844), .Y(n5695) );
  INVX1 U4355 ( .A(n5694), .Y(n5635) );
  INVX1 U4356 ( .A(n5694), .Y(n5636) );
  INVX1 U4357 ( .A(n5694), .Y(n5637) );
  INVX1 U4358 ( .A(n5843), .Y(n5704) );
  INVX1 U4359 ( .A(n5843), .Y(n5703) );
  INVX1 U4360 ( .A(n5843), .Y(n5702) );
  INVX1 U4361 ( .A(n5843), .Y(n5701) );
  INVX1 U4362 ( .A(n5843), .Y(n5700) );
  INVX1 U4363 ( .A(n5843), .Y(n5699) );
  INVX1 U4364 ( .A(n5843), .Y(n5698) );
  INVX1 U4365 ( .A(n5843), .Y(n5697) );
  INVX1 U4366 ( .A(n5843), .Y(n5696) );
  AND2X1 U4367 ( .A(n1642), .B(n1575), .Y(n1578) );
  INVX1 U4368 ( .A(n5775), .Y(n5774) );
  INVX1 U4369 ( .A(n661), .Y(n5816) );
  INVX1 U4370 ( .A(n747), .Y(n5812) );
  INVX1 U4371 ( .A(n790), .Y(n5810) );
  INVX1 U4372 ( .A(n833), .Y(n5808) );
  INVX1 U4373 ( .A(n1006), .Y(n5800) );
  INVX1 U4374 ( .A(n1092), .Y(n5796) );
  INVX1 U4375 ( .A(n1135), .Y(n5794) );
  INVX1 U4376 ( .A(n1178), .Y(n5792) );
  INVX1 U4377 ( .A(n531), .Y(n5822) );
  INVX1 U4378 ( .A(n575), .Y(n5820) );
  INVX1 U4379 ( .A(n876), .Y(n5806) );
  INVX1 U4380 ( .A(n920), .Y(n5804) );
  INVX1 U4381 ( .A(n618), .Y(n5818) );
  INVX1 U4382 ( .A(n704), .Y(n5814) );
  INVX1 U4383 ( .A(n963), .Y(n5802) );
  INVX1 U4384 ( .A(n1049), .Y(n5798) );
  INVX1 U4385 ( .A(n223), .Y(n5836) );
  INVX1 U4386 ( .A(n267), .Y(n5834) );
  INVX1 U4387 ( .A(n311), .Y(n5832) );
  INVX1 U4388 ( .A(n355), .Y(n5830) );
  INVX1 U4389 ( .A(n399), .Y(n5828) );
  INVX1 U4390 ( .A(n443), .Y(n5826) );
  INVX1 U4391 ( .A(n487), .Y(n5824) );
  INVX1 U4392 ( .A(n661), .Y(n5817) );
  INVX1 U4393 ( .A(n747), .Y(n5813) );
  INVX1 U4394 ( .A(n790), .Y(n5811) );
  INVX1 U4395 ( .A(n833), .Y(n5809) );
  INVX1 U4396 ( .A(n1006), .Y(n5801) );
  INVX1 U4397 ( .A(n1092), .Y(n5797) );
  INVX1 U4398 ( .A(n1135), .Y(n5795) );
  INVX1 U4399 ( .A(n1178), .Y(n5793) );
  INVX1 U4400 ( .A(n1351), .Y(n5784) );
  INVX1 U4401 ( .A(n1437), .Y(n5780) );
  INVX1 U4402 ( .A(n1480), .Y(n5778) );
  INVX1 U4403 ( .A(n531), .Y(n5823) );
  INVX1 U4404 ( .A(n575), .Y(n5821) );
  INVX1 U4405 ( .A(n876), .Y(n5807) );
  INVX1 U4406 ( .A(n920), .Y(n5805) );
  INVX1 U4407 ( .A(n618), .Y(n5819) );
  INVX1 U4408 ( .A(n704), .Y(n5815) );
  INVX1 U4409 ( .A(n963), .Y(n5803) );
  INVX1 U4410 ( .A(n1049), .Y(n5799) );
  INVX1 U4411 ( .A(n1308), .Y(n5786) );
  INVX1 U4412 ( .A(n1394), .Y(n5782) );
  INVX1 U4413 ( .A(n223), .Y(n5837) );
  INVX1 U4414 ( .A(n267), .Y(n5835) );
  INVX1 U4415 ( .A(n311), .Y(n5833) );
  INVX1 U4416 ( .A(n355), .Y(n5831) );
  INVX1 U4417 ( .A(n399), .Y(n5829) );
  INVX1 U4418 ( .A(n443), .Y(n5827) );
  INVX1 U4419 ( .A(n487), .Y(n5825) );
  INVX1 U4420 ( .A(n1221), .Y(n5790) );
  INVX1 U4421 ( .A(n1265), .Y(n5788) );
  INVX1 U4422 ( .A(n178), .Y(n5838) );
  INVX1 U4423 ( .A(n1351), .Y(n5785) );
  INVX1 U4424 ( .A(n1437), .Y(n5781) );
  INVX1 U4425 ( .A(n1480), .Y(n5779) );
  INVX1 U4426 ( .A(n1221), .Y(n5791) );
  INVX1 U4427 ( .A(n1265), .Y(n5789) );
  INVX1 U4428 ( .A(n1308), .Y(n5787) );
  INVX1 U4429 ( .A(n1394), .Y(n5783) );
  INVX1 U4430 ( .A(n178), .Y(n5839) );
  INVX1 U4431 ( .A(n5843), .Y(n5723) );
  AND2X1 U4432 ( .A(n1643), .B(n1575), .Y(n1577) );
  INVX1 U4433 ( .A(n4323), .Y(n5775) );
  AND2X1 U4434 ( .A(n1647), .B(n5845), .Y(n1642) );
  INVX1 U4435 ( .A(reset), .Y(n5845) );
  INVX1 U4436 ( .A(data_in[8]), .Y(n5738) );
  INVX1 U4437 ( .A(data_in[2]), .Y(n5744) );
  INVX1 U4438 ( .A(data_in[3]), .Y(n5743) );
  INVX1 U4439 ( .A(data_in[4]), .Y(n5742) );
  INVX1 U4440 ( .A(data_in[5]), .Y(n5741) );
  INVX1 U4441 ( .A(data_in[9]), .Y(n5737) );
  INVX1 U4442 ( .A(data_in[10]), .Y(n5736) );
  INVX1 U4443 ( .A(data_in[11]), .Y(n5735) );
  INVX1 U4444 ( .A(data_in[12]), .Y(n5734) );
  INVX1 U4445 ( .A(data_in[13]), .Y(n5733) );
  INVX1 U4446 ( .A(data_in[6]), .Y(n5740) );
  INVX1 U4447 ( .A(data_in[14]), .Y(n5732) );
  INVX1 U4448 ( .A(data_in[1]), .Y(n5745) );
  INVX1 U4449 ( .A(data_in[7]), .Y(n5739) );
  INVX1 U4450 ( .A(data_in[15]), .Y(n5731) );
  INVX1 U4451 ( .A(data_in[0]), .Y(n5746) );
  INVX1 U4452 ( .A(n4321), .Y(n5894) );
  INVX1 U4453 ( .A(data_in[16]), .Y(n5749) );
  INVX1 U4454 ( .A(data_in[17]), .Y(n5750) );
  INVX1 U4455 ( .A(data_in[18]), .Y(n5751) );
  INVX1 U4456 ( .A(data_in[19]), .Y(n5752) );
  INVX1 U4457 ( .A(data_in[20]), .Y(n5753) );
  INVX1 U4458 ( .A(data_in[21]), .Y(n5754) );
  INVX1 U4459 ( .A(data_in[22]), .Y(n5755) );
  INVX1 U4460 ( .A(data_in[23]), .Y(n5756) );
  INVX1 U4461 ( .A(data_in[24]), .Y(n5757) );
  INVX1 U4462 ( .A(data_in[25]), .Y(n5758) );
  INVX1 U4463 ( .A(data_in[26]), .Y(n5759) );
  INVX1 U4464 ( .A(data_in[27]), .Y(n5760) );
  INVX1 U4465 ( .A(data_in[28]), .Y(n5761) );
  INVX1 U4466 ( .A(data_in[29]), .Y(n5762) );
  INVX1 U4467 ( .A(data_in[30]), .Y(n5763) );
  INVX1 U4468 ( .A(data_in[31]), .Y(n5764) );
  INVX1 U4469 ( .A(data_in[32]), .Y(n5765) );
  INVX1 U4470 ( .A(data_in[33]), .Y(n5766) );
  INVX1 U4471 ( .A(data_in[34]), .Y(n5767) );
  INVX1 U4472 ( .A(data_in[35]), .Y(n5768) );
  INVX1 U4473 ( .A(data_in[36]), .Y(n5769) );
  INVX1 U4474 ( .A(data_in[37]), .Y(n5770) );
  INVX1 U4475 ( .A(data_in[38]), .Y(n5771) );
  INVX1 U4476 ( .A(data_in[39]), .Y(n5772) );
  INVX1 U4477 ( .A(data_in[40]), .Y(n5748) );
  INVX1 U4478 ( .A(data_in[41]), .Y(n5747) );
  INVX1 U4479 ( .A(n102), .Y(n5893) );
  INVX1 U4480 ( .A(n5625), .Y(n24) );
  INVX1 U4481 ( .A(n101), .Y(n5892) );
  INVX1 U4482 ( .A(n5624), .Y(n25) );
  INVX1 U4483 ( .A(n100), .Y(n5891) );
  INVX1 U4484 ( .A(n5623), .Y(n26) );
  INVX1 U4485 ( .A(n99), .Y(n5890) );
  INVX1 U4486 ( .A(n5622), .Y(n27) );
  INVX1 U4487 ( .A(n98), .Y(n5889) );
  INVX1 U4488 ( .A(n5621), .Y(n28) );
  INVX1 U4489 ( .A(n97), .Y(n5888) );
  INVX1 U4490 ( .A(n5620), .Y(n29) );
  INVX1 U4491 ( .A(n91), .Y(n5887) );
  INVX1 U4492 ( .A(n5619), .Y(n30) );
  INVX1 U4493 ( .A(n90), .Y(n5886) );
  INVX1 U4494 ( .A(n5618), .Y(n31) );
  INVX1 U4495 ( .A(n89), .Y(n5885) );
  INVX1 U4496 ( .A(n5617), .Y(n32) );
  INVX1 U4497 ( .A(n88), .Y(n5884) );
  INVX1 U4498 ( .A(n5616), .Y(n33) );
  INVX1 U4499 ( .A(n87), .Y(n5883) );
  INVX1 U4500 ( .A(n5615), .Y(n34) );
  INVX1 U4501 ( .A(n86), .Y(n5882) );
  INVX1 U4502 ( .A(n5614), .Y(n35) );
  INVX1 U4503 ( .A(n85), .Y(n5881) );
  INVX1 U4504 ( .A(n5613), .Y(n36) );
  INVX1 U4505 ( .A(n80), .Y(n5880) );
  INVX1 U4506 ( .A(n5612), .Y(n37) );
  INVX1 U4507 ( .A(n75), .Y(n5879) );
  INVX1 U4508 ( .A(n5611), .Y(n38) );
  INVX1 U4509 ( .A(n74), .Y(n5878) );
  INVX1 U4510 ( .A(n5610), .Y(n39) );
  INVX1 U4511 ( .A(n73), .Y(n5877) );
  INVX1 U4512 ( .A(n5609), .Y(n40) );
  INVX1 U4513 ( .A(n72), .Y(n5876) );
  INVX1 U4514 ( .A(n5608), .Y(n41) );
  INVX1 U4515 ( .A(n71), .Y(n5875) );
  INVX1 U4516 ( .A(n5607), .Y(n42) );
  INVX1 U4517 ( .A(n70), .Y(n5874) );
  INVX1 U4518 ( .A(n5606), .Y(n43) );
  INVX1 U4519 ( .A(n69), .Y(n5873) );
  INVX1 U4520 ( .A(n5605), .Y(n44) );
  INVX1 U4521 ( .A(n68), .Y(n5872) );
  INVX1 U4522 ( .A(n5604), .Y(n45) );
  INVX1 U4523 ( .A(n67), .Y(n5871) );
  INVX1 U4524 ( .A(n5603), .Y(n46) );
  INVX1 U4525 ( .A(n66), .Y(n5870) );
  INVX1 U4526 ( .A(n5602), .Y(n47) );
  INVX1 U4527 ( .A(n18), .Y(n5869) );
  INVX1 U4528 ( .A(n5601), .Y(n48) );
  INVX1 U4529 ( .A(n17), .Y(n5868) );
  INVX1 U4530 ( .A(n5600), .Y(n49) );
  INVX1 U4531 ( .A(n16), .Y(n5867) );
  INVX1 U4532 ( .A(n5599), .Y(n50) );
  INVX1 U4533 ( .A(n15), .Y(n5866) );
  INVX1 U4534 ( .A(n5598), .Y(n51) );
  INVX1 U4535 ( .A(n14), .Y(n5865) );
  INVX1 U4536 ( .A(n5597), .Y(n52) );
  INVX1 U4537 ( .A(n13), .Y(n5864) );
  INVX1 U4538 ( .A(n5596), .Y(n53) );
  INVX1 U4539 ( .A(n12), .Y(n5863) );
  INVX1 U4540 ( .A(n5595), .Y(n54) );
  INVX1 U4541 ( .A(n11), .Y(n5862) );
  INVX1 U4542 ( .A(n5594), .Y(n55) );
  INVX1 U4543 ( .A(n10), .Y(n5861) );
  INVX1 U4544 ( .A(n5593), .Y(n56) );
  INVX1 U4545 ( .A(n9), .Y(n5860) );
  INVX1 U4546 ( .A(n5592), .Y(n57) );
  INVX1 U4547 ( .A(n8), .Y(n5859) );
  INVX1 U4548 ( .A(n5591), .Y(n58) );
  INVX1 U4549 ( .A(n7), .Y(n5858) );
  INVX1 U4550 ( .A(n5590), .Y(n59) );
  INVX1 U4551 ( .A(n6), .Y(n5857) );
  INVX1 U4552 ( .A(n5589), .Y(n60) );
  INVX1 U4553 ( .A(n5), .Y(n5856) );
  INVX1 U4554 ( .A(n5588), .Y(n61) );
  INVX1 U4555 ( .A(n4), .Y(n5855) );
  INVX1 U4556 ( .A(n5587), .Y(n62) );
  INVX1 U4557 ( .A(n3), .Y(n5854) );
  INVX1 U4558 ( .A(n5586), .Y(n63) );
  INVX1 U4559 ( .A(n2), .Y(n5853) );
  INVX1 U4560 ( .A(n5585), .Y(n64) );
  INVX1 U4561 ( .A(n1), .Y(n5852) );
  INVX1 U4562 ( .A(n5584), .Y(n65) );
  INVX1 U4563 ( .A(empty), .Y(n5897) );
  INVX1 U4564 ( .A(n19), .Y(n5844) );
  INVX1 U4565 ( .A(full), .Y(n5895) );
  INVX1 U4566 ( .A(wr_ptr[2]), .Y(n5900) );
  INVX1 U4567 ( .A(wr_ptr[0]), .Y(n5898) );
  INVX1 U4568 ( .A(wr_ptr[1]), .Y(n5899) );
  INVX1 U4569 ( .A(wr_ptr[4]), .Y(n5902) );
  INVX1 U4570 ( .A(wr_ptr[3]), .Y(n5901) );
  INVX1 U4571 ( .A(fillcount[4]), .Y(n5903) );
  INVX1 U4572 ( .A(fillcount[0]), .Y(n103) );
  INVX1 U4573 ( .A(fillcount[5]), .Y(n5896) );
  INVX1 U4574 ( .A(fillcount[2]), .Y(n5851) );
  INVX1 U4575 ( .A(fillcount[3]), .Y(n5850) );
  INVX1 U4576 ( .A(fillcount[1]), .Y(n5904) );
  INVX1 U4577 ( .A(n20), .Y(n5843) );
  INVX1 U4578 ( .A(n21), .Y(n5842) );
  INVX1 U4579 ( .A(n22), .Y(n5841) );
  INVX1 U4580 ( .A(n23), .Y(n5840) );
  AND2X1 U4581 ( .A(n5904), .B(fillcount[0]), .Y(n1638) );
  MUX2X1 U4582 ( .B(n4325), .A(n4326), .S(n5696), .Y(n4324) );
  MUX2X1 U4583 ( .B(n4328), .A(n4329), .S(n5696), .Y(n4327) );
  MUX2X1 U4584 ( .B(n4331), .A(n4332), .S(n5696), .Y(n4330) );
  MUX2X1 U4585 ( .B(n4334), .A(n4335), .S(n5696), .Y(n4333) );
  MUX2X1 U4586 ( .B(n4337), .A(n4338), .S(n22), .Y(n4336) );
  MUX2X1 U4587 ( .B(n4340), .A(n4341), .S(n5696), .Y(n4339) );
  MUX2X1 U4588 ( .B(n4343), .A(n4344), .S(n5696), .Y(n4342) );
  MUX2X1 U4589 ( .B(n4346), .A(n4347), .S(n5696), .Y(n4345) );
  MUX2X1 U4590 ( .B(n4349), .A(n4350), .S(n5696), .Y(n4348) );
  MUX2X1 U4591 ( .B(n4352), .A(n4353), .S(n22), .Y(n4351) );
  MUX2X1 U4592 ( .B(n4355), .A(n4356), .S(n5696), .Y(n4354) );
  MUX2X1 U4593 ( .B(n4358), .A(n4359), .S(n5696), .Y(n4357) );
  MUX2X1 U4594 ( .B(n4361), .A(n4362), .S(n5696), .Y(n4360) );
  MUX2X1 U4595 ( .B(n4364), .A(n4365), .S(n5696), .Y(n4363) );
  MUX2X1 U4596 ( .B(n4367), .A(n4368), .S(n22), .Y(n4366) );
  MUX2X1 U4597 ( .B(n4370), .A(n4371), .S(n5697), .Y(n4369) );
  MUX2X1 U4598 ( .B(n4373), .A(n4374), .S(n5697), .Y(n4372) );
  MUX2X1 U4599 ( .B(n4376), .A(n4377), .S(n5697), .Y(n4375) );
  MUX2X1 U4600 ( .B(n4379), .A(n4380), .S(n5697), .Y(n4378) );
  MUX2X1 U4601 ( .B(n4382), .A(n4383), .S(n22), .Y(n4381) );
  MUX2X1 U4602 ( .B(n4385), .A(n4386), .S(n5697), .Y(n4384) );
  MUX2X1 U4603 ( .B(n4388), .A(n4389), .S(n5697), .Y(n4387) );
  MUX2X1 U4604 ( .B(n4391), .A(n4392), .S(n5697), .Y(n4390) );
  MUX2X1 U4605 ( .B(n4394), .A(n4395), .S(n5697), .Y(n4393) );
  MUX2X1 U4606 ( .B(n4397), .A(n4398), .S(n22), .Y(n4396) );
  MUX2X1 U4607 ( .B(n4400), .A(n4401), .S(n5697), .Y(n4399) );
  MUX2X1 U4608 ( .B(n4403), .A(n4404), .S(n5697), .Y(n4402) );
  MUX2X1 U4609 ( .B(n4406), .A(n4407), .S(n5697), .Y(n4405) );
  MUX2X1 U4610 ( .B(n4409), .A(n4410), .S(n5697), .Y(n4408) );
  MUX2X1 U4611 ( .B(n4412), .A(n4413), .S(n22), .Y(n4411) );
  MUX2X1 U4612 ( .B(n4415), .A(n4416), .S(n5698), .Y(n4414) );
  MUX2X1 U4613 ( .B(n4418), .A(n4419), .S(n5698), .Y(n4417) );
  MUX2X1 U4614 ( .B(n4421), .A(n4422), .S(n5698), .Y(n4420) );
  MUX2X1 U4615 ( .B(n4424), .A(n4425), .S(n5698), .Y(n4423) );
  MUX2X1 U4616 ( .B(n4427), .A(n4428), .S(n22), .Y(n4426) );
  MUX2X1 U4617 ( .B(n4430), .A(n4431), .S(n5698), .Y(n4429) );
  MUX2X1 U4618 ( .B(n4433), .A(n4434), .S(n5698), .Y(n4432) );
  MUX2X1 U4619 ( .B(n4436), .A(n4437), .S(n5698), .Y(n4435) );
  MUX2X1 U4620 ( .B(n4439), .A(n4440), .S(n5698), .Y(n4438) );
  MUX2X1 U4621 ( .B(n4442), .A(n4443), .S(n22), .Y(n4441) );
  MUX2X1 U4622 ( .B(n4445), .A(n4446), .S(n5698), .Y(n4444) );
  MUX2X1 U4623 ( .B(n4448), .A(n4449), .S(n5698), .Y(n4447) );
  MUX2X1 U4624 ( .B(n4451), .A(n4452), .S(n5698), .Y(n4450) );
  MUX2X1 U4625 ( .B(n4454), .A(n4455), .S(n5698), .Y(n4453) );
  MUX2X1 U4626 ( .B(n4457), .A(n4458), .S(n22), .Y(n4456) );
  MUX2X1 U4627 ( .B(n4460), .A(n4461), .S(n5699), .Y(n4459) );
  MUX2X1 U4628 ( .B(n4463), .A(n4464), .S(n5699), .Y(n4462) );
  MUX2X1 U4629 ( .B(n4466), .A(n4467), .S(n5699), .Y(n4465) );
  MUX2X1 U4630 ( .B(n4469), .A(n4470), .S(n5699), .Y(n4468) );
  MUX2X1 U4631 ( .B(n4472), .A(n4473), .S(n22), .Y(n4471) );
  MUX2X1 U4632 ( .B(n4475), .A(n4476), .S(n5699), .Y(n4474) );
  MUX2X1 U4633 ( .B(n4478), .A(n4479), .S(n5699), .Y(n4477) );
  MUX2X1 U4634 ( .B(n4481), .A(n4482), .S(n5699), .Y(n4480) );
  MUX2X1 U4635 ( .B(n4484), .A(n4485), .S(n5699), .Y(n4483) );
  MUX2X1 U4636 ( .B(n4487), .A(n4488), .S(n22), .Y(n4486) );
  MUX2X1 U4637 ( .B(n4490), .A(n4491), .S(n5699), .Y(n4489) );
  MUX2X1 U4638 ( .B(n4493), .A(n4494), .S(n5699), .Y(n4492) );
  MUX2X1 U4639 ( .B(n4496), .A(n4497), .S(n5699), .Y(n4495) );
  MUX2X1 U4640 ( .B(n4499), .A(n4500), .S(n5699), .Y(n4498) );
  MUX2X1 U4641 ( .B(n4502), .A(n4503), .S(n22), .Y(n4501) );
  MUX2X1 U4642 ( .B(n4505), .A(n4506), .S(n5700), .Y(n4504) );
  MUX2X1 U4643 ( .B(n4508), .A(n4509), .S(n5700), .Y(n4507) );
  MUX2X1 U4644 ( .B(n4511), .A(n4512), .S(n5700), .Y(n4510) );
  MUX2X1 U4645 ( .B(n4514), .A(n4515), .S(n5700), .Y(n4513) );
  MUX2X1 U4646 ( .B(n4517), .A(n4518), .S(n22), .Y(n4516) );
  MUX2X1 U4647 ( .B(n4520), .A(n4521), .S(n5700), .Y(n4519) );
  MUX2X1 U4648 ( .B(n4523), .A(n4524), .S(n5700), .Y(n4522) );
  MUX2X1 U4649 ( .B(n4526), .A(n4527), .S(n5700), .Y(n4525) );
  MUX2X1 U4650 ( .B(n4529), .A(n4530), .S(n5700), .Y(n4528) );
  MUX2X1 U4651 ( .B(n4532), .A(n4533), .S(n22), .Y(n4531) );
  MUX2X1 U4652 ( .B(n4535), .A(n4536), .S(n5700), .Y(n4534) );
  MUX2X1 U4653 ( .B(n4538), .A(n4539), .S(n5700), .Y(n4537) );
  MUX2X1 U4654 ( .B(n4541), .A(n4542), .S(n5700), .Y(n4540) );
  MUX2X1 U4655 ( .B(n4544), .A(n4545), .S(n5700), .Y(n4543) );
  MUX2X1 U4656 ( .B(n4547), .A(n4548), .S(n22), .Y(n4546) );
  MUX2X1 U4657 ( .B(n4550), .A(n4551), .S(n5701), .Y(n4549) );
  MUX2X1 U4658 ( .B(n4553), .A(n4554), .S(n5701), .Y(n4552) );
  MUX2X1 U4659 ( .B(n4556), .A(n4557), .S(n5701), .Y(n4555) );
  MUX2X1 U4660 ( .B(n4559), .A(n4560), .S(n5701), .Y(n4558) );
  MUX2X1 U4661 ( .B(n4562), .A(n4563), .S(n22), .Y(n4561) );
  MUX2X1 U4662 ( .B(n4565), .A(n4566), .S(n5701), .Y(n4564) );
  MUX2X1 U4663 ( .B(n4568), .A(n4569), .S(n5701), .Y(n4567) );
  MUX2X1 U4664 ( .B(n4571), .A(n4572), .S(n5701), .Y(n4570) );
  MUX2X1 U4665 ( .B(n4574), .A(n4575), .S(n5701), .Y(n4573) );
  MUX2X1 U4666 ( .B(n4577), .A(n4578), .S(n22), .Y(n4576) );
  MUX2X1 U4667 ( .B(n4580), .A(n4581), .S(n5701), .Y(n4579) );
  MUX2X1 U4668 ( .B(n4583), .A(n4584), .S(n5701), .Y(n4582) );
  MUX2X1 U4669 ( .B(n4586), .A(n4587), .S(n5701), .Y(n4585) );
  MUX2X1 U4670 ( .B(n4589), .A(n4590), .S(n5701), .Y(n4588) );
  MUX2X1 U4671 ( .B(n4592), .A(n4593), .S(n22), .Y(n4591) );
  MUX2X1 U4672 ( .B(n4595), .A(n4596), .S(n5702), .Y(n4594) );
  MUX2X1 U4673 ( .B(n4598), .A(n4599), .S(n5702), .Y(n4597) );
  MUX2X1 U4674 ( .B(n4601), .A(n4602), .S(n5702), .Y(n4600) );
  MUX2X1 U4675 ( .B(n4604), .A(n4605), .S(n5702), .Y(n4603) );
  MUX2X1 U4676 ( .B(n4607), .A(n4608), .S(n22), .Y(n4606) );
  MUX2X1 U4677 ( .B(n4610), .A(n4611), .S(n5702), .Y(n4609) );
  MUX2X1 U4678 ( .B(n4613), .A(n4614), .S(n5702), .Y(n4612) );
  MUX2X1 U4679 ( .B(n4616), .A(n4617), .S(n5702), .Y(n4615) );
  MUX2X1 U4680 ( .B(n4619), .A(n4620), .S(n5702), .Y(n4618) );
  MUX2X1 U4681 ( .B(n4622), .A(n4623), .S(n22), .Y(n4621) );
  MUX2X1 U4682 ( .B(n4625), .A(n4626), .S(n5702), .Y(n4624) );
  MUX2X1 U4683 ( .B(n4628), .A(n4629), .S(n5702), .Y(n4627) );
  MUX2X1 U4684 ( .B(n4631), .A(n4632), .S(n5702), .Y(n4630) );
  MUX2X1 U4685 ( .B(n4634), .A(n4635), .S(n5702), .Y(n4633) );
  MUX2X1 U4686 ( .B(n4637), .A(n4638), .S(n22), .Y(n4636) );
  MUX2X1 U4687 ( .B(n4640), .A(n4641), .S(n5703), .Y(n4639) );
  MUX2X1 U4688 ( .B(n4643), .A(n4644), .S(n5703), .Y(n4642) );
  MUX2X1 U4689 ( .B(n4646), .A(n4647), .S(n5703), .Y(n4645) );
  MUX2X1 U4690 ( .B(n4649), .A(n4650), .S(n5703), .Y(n4648) );
  MUX2X1 U4691 ( .B(n4652), .A(n4653), .S(n22), .Y(n4651) );
  MUX2X1 U4692 ( .B(n4655), .A(n4656), .S(n5703), .Y(n4654) );
  MUX2X1 U4693 ( .B(n4658), .A(n4659), .S(n5703), .Y(n4657) );
  MUX2X1 U4694 ( .B(n4661), .A(n4662), .S(n5703), .Y(n4660) );
  MUX2X1 U4695 ( .B(n4664), .A(n4665), .S(n5703), .Y(n4663) );
  MUX2X1 U4696 ( .B(n4667), .A(n4668), .S(n22), .Y(n4666) );
  MUX2X1 U4697 ( .B(n4670), .A(n4671), .S(n5703), .Y(n4669) );
  MUX2X1 U4698 ( .B(n4673), .A(n4674), .S(n5703), .Y(n4672) );
  MUX2X1 U4699 ( .B(n4676), .A(n4677), .S(n5703), .Y(n4675) );
  MUX2X1 U4700 ( .B(n4679), .A(n4680), .S(n5703), .Y(n4678) );
  MUX2X1 U4701 ( .B(n4682), .A(n4683), .S(n22), .Y(n4681) );
  MUX2X1 U4702 ( .B(n4685), .A(n4686), .S(n5704), .Y(n4684) );
  MUX2X1 U4703 ( .B(n4688), .A(n4689), .S(n5704), .Y(n4687) );
  MUX2X1 U4704 ( .B(n4691), .A(n4692), .S(n5704), .Y(n4690) );
  MUX2X1 U4705 ( .B(n4694), .A(n4695), .S(n5704), .Y(n4693) );
  MUX2X1 U4706 ( .B(n4697), .A(n4698), .S(n22), .Y(n4696) );
  MUX2X1 U4707 ( .B(n4700), .A(n4701), .S(n5704), .Y(n4699) );
  MUX2X1 U4708 ( .B(n4703), .A(n4704), .S(n5704), .Y(n4702) );
  MUX2X1 U4709 ( .B(n4706), .A(n4707), .S(n5704), .Y(n4705) );
  MUX2X1 U4710 ( .B(n4709), .A(n4710), .S(n5704), .Y(n4708) );
  MUX2X1 U4711 ( .B(n4712), .A(n4713), .S(n22), .Y(n4711) );
  MUX2X1 U4712 ( .B(n4715), .A(n4716), .S(n5704), .Y(n4714) );
  MUX2X1 U4713 ( .B(n4718), .A(n4719), .S(n5704), .Y(n4717) );
  MUX2X1 U4714 ( .B(n4721), .A(n4722), .S(n5704), .Y(n4720) );
  MUX2X1 U4715 ( .B(n4724), .A(n4725), .S(n5704), .Y(n4723) );
  MUX2X1 U4716 ( .B(n4727), .A(n4728), .S(n22), .Y(n4726) );
  MUX2X1 U4717 ( .B(n4730), .A(n4731), .S(n5705), .Y(n4729) );
  MUX2X1 U4718 ( .B(n4733), .A(n4734), .S(n5705), .Y(n4732) );
  MUX2X1 U4719 ( .B(n4736), .A(n4737), .S(n5705), .Y(n4735) );
  MUX2X1 U4720 ( .B(n4739), .A(n4740), .S(n5705), .Y(n4738) );
  MUX2X1 U4721 ( .B(n4742), .A(n4743), .S(n22), .Y(n4741) );
  MUX2X1 U4722 ( .B(n4745), .A(n4746), .S(n5705), .Y(n4744) );
  MUX2X1 U4723 ( .B(n4748), .A(n4749), .S(n5705), .Y(n4747) );
  MUX2X1 U4724 ( .B(n4751), .A(n4752), .S(n5705), .Y(n4750) );
  MUX2X1 U4725 ( .B(n4754), .A(n4755), .S(n5705), .Y(n4753) );
  MUX2X1 U4726 ( .B(n4757), .A(n4758), .S(n22), .Y(n4756) );
  MUX2X1 U4727 ( .B(n4760), .A(n4761), .S(n5705), .Y(n4759) );
  MUX2X1 U4728 ( .B(n4763), .A(n4764), .S(n5705), .Y(n4762) );
  MUX2X1 U4729 ( .B(n4766), .A(n4767), .S(n5705), .Y(n4765) );
  MUX2X1 U4730 ( .B(n4769), .A(n4770), .S(n5705), .Y(n4768) );
  MUX2X1 U4731 ( .B(n4772), .A(n4773), .S(n22), .Y(n4771) );
  MUX2X1 U4732 ( .B(n4775), .A(n4776), .S(n5706), .Y(n4774) );
  MUX2X1 U4733 ( .B(n4778), .A(n4779), .S(n5706), .Y(n4777) );
  MUX2X1 U4734 ( .B(n4781), .A(n4782), .S(n5706), .Y(n4780) );
  MUX2X1 U4735 ( .B(n4784), .A(n4785), .S(n5706), .Y(n4783) );
  MUX2X1 U4736 ( .B(n4787), .A(n4788), .S(n22), .Y(n4786) );
  MUX2X1 U4737 ( .B(n4790), .A(n4791), .S(n5706), .Y(n4789) );
  MUX2X1 U4738 ( .B(n4793), .A(n4794), .S(n5706), .Y(n4792) );
  MUX2X1 U4739 ( .B(n4796), .A(n4797), .S(n5706), .Y(n4795) );
  MUX2X1 U4740 ( .B(n4799), .A(n4800), .S(n5706), .Y(n4798) );
  MUX2X1 U4741 ( .B(n4802), .A(n4803), .S(n22), .Y(n4801) );
  MUX2X1 U4742 ( .B(n4805), .A(n4806), .S(n5706), .Y(n4804) );
  MUX2X1 U4743 ( .B(n4808), .A(n4809), .S(n5706), .Y(n4807) );
  MUX2X1 U4744 ( .B(n4811), .A(n4812), .S(n5706), .Y(n4810) );
  MUX2X1 U4745 ( .B(n4814), .A(n4815), .S(n5706), .Y(n4813) );
  MUX2X1 U4746 ( .B(n4817), .A(n4818), .S(n22), .Y(n4816) );
  MUX2X1 U4747 ( .B(n4820), .A(n4821), .S(n5707), .Y(n4819) );
  MUX2X1 U4748 ( .B(n4823), .A(n4824), .S(n5707), .Y(n4822) );
  MUX2X1 U4749 ( .B(n4826), .A(n4827), .S(n5707), .Y(n4825) );
  MUX2X1 U4750 ( .B(n4829), .A(n4830), .S(n5707), .Y(n4828) );
  MUX2X1 U4751 ( .B(n4832), .A(n4833), .S(n22), .Y(n4831) );
  MUX2X1 U4752 ( .B(n4835), .A(n4836), .S(n5707), .Y(n4834) );
  MUX2X1 U4753 ( .B(n4838), .A(n4839), .S(n5707), .Y(n4837) );
  MUX2X1 U4754 ( .B(n4841), .A(n4842), .S(n5707), .Y(n4840) );
  MUX2X1 U4755 ( .B(n4844), .A(n4845), .S(n5707), .Y(n4843) );
  MUX2X1 U4756 ( .B(n4847), .A(n4848), .S(n22), .Y(n4846) );
  MUX2X1 U4757 ( .B(n4850), .A(n4851), .S(n5707), .Y(n4849) );
  MUX2X1 U4758 ( .B(n4853), .A(n4854), .S(n5707), .Y(n4852) );
  MUX2X1 U4759 ( .B(n4856), .A(n4857), .S(n5707), .Y(n4855) );
  MUX2X1 U4760 ( .B(n4859), .A(n4860), .S(n5707), .Y(n4858) );
  MUX2X1 U4761 ( .B(n4862), .A(n4863), .S(n22), .Y(n4861) );
  MUX2X1 U4762 ( .B(n4865), .A(n4866), .S(n5708), .Y(n4864) );
  MUX2X1 U4763 ( .B(n4868), .A(n4869), .S(n5708), .Y(n4867) );
  MUX2X1 U4764 ( .B(n4871), .A(n4872), .S(n5708), .Y(n4870) );
  MUX2X1 U4765 ( .B(n4874), .A(n4875), .S(n5708), .Y(n4873) );
  MUX2X1 U4766 ( .B(n4877), .A(n4878), .S(n22), .Y(n4876) );
  MUX2X1 U4767 ( .B(n4880), .A(n4881), .S(n5708), .Y(n4879) );
  MUX2X1 U4768 ( .B(n4883), .A(n4884), .S(n5708), .Y(n4882) );
  MUX2X1 U4769 ( .B(n4886), .A(n4887), .S(n5708), .Y(n4885) );
  MUX2X1 U4770 ( .B(n4889), .A(n4890), .S(n5708), .Y(n4888) );
  MUX2X1 U4771 ( .B(n4892), .A(n4893), .S(n22), .Y(n4891) );
  MUX2X1 U4772 ( .B(n4895), .A(n4896), .S(n5708), .Y(n4894) );
  MUX2X1 U4773 ( .B(n4898), .A(n4899), .S(n5708), .Y(n4897) );
  MUX2X1 U4774 ( .B(n4901), .A(n4902), .S(n5708), .Y(n4900) );
  MUX2X1 U4775 ( .B(n4904), .A(n4905), .S(n5708), .Y(n4903) );
  MUX2X1 U4776 ( .B(n4907), .A(n4908), .S(n22), .Y(n4906) );
  MUX2X1 U4777 ( .B(n4910), .A(n4911), .S(n5709), .Y(n4909) );
  MUX2X1 U4778 ( .B(n4913), .A(n4914), .S(n5709), .Y(n4912) );
  MUX2X1 U4779 ( .B(n4916), .A(n4917), .S(n5709), .Y(n4915) );
  MUX2X1 U4780 ( .B(n4919), .A(n4920), .S(n5709), .Y(n4918) );
  MUX2X1 U4781 ( .B(n4922), .A(n4923), .S(n22), .Y(n4921) );
  MUX2X1 U4782 ( .B(n4925), .A(n4926), .S(n5709), .Y(n4924) );
  MUX2X1 U4783 ( .B(n4928), .A(n4929), .S(n5709), .Y(n4927) );
  MUX2X1 U4784 ( .B(n4931), .A(n4932), .S(n5709), .Y(n4930) );
  MUX2X1 U4785 ( .B(n4934), .A(n4935), .S(n5709), .Y(n4933) );
  MUX2X1 U4786 ( .B(n4937), .A(n4938), .S(n22), .Y(n4936) );
  MUX2X1 U4787 ( .B(n4940), .A(n4941), .S(n5709), .Y(n4939) );
  MUX2X1 U4788 ( .B(n4943), .A(n4944), .S(n5709), .Y(n4942) );
  MUX2X1 U4789 ( .B(n4946), .A(n4947), .S(n5709), .Y(n4945) );
  MUX2X1 U4790 ( .B(n4949), .A(n4950), .S(n5709), .Y(n4948) );
  MUX2X1 U4791 ( .B(n4952), .A(n4953), .S(n22), .Y(n4951) );
  MUX2X1 U4792 ( .B(n4955), .A(n4956), .S(n5710), .Y(n4954) );
  MUX2X1 U4793 ( .B(n4958), .A(n4959), .S(n5710), .Y(n4957) );
  MUX2X1 U4794 ( .B(n4961), .A(n4962), .S(n5710), .Y(n4960) );
  MUX2X1 U4795 ( .B(n4964), .A(n4965), .S(n5710), .Y(n4963) );
  MUX2X1 U4796 ( .B(n4967), .A(n4968), .S(n22), .Y(n4966) );
  MUX2X1 U4797 ( .B(n4970), .A(n4971), .S(n5710), .Y(n4969) );
  MUX2X1 U4798 ( .B(n4973), .A(n4974), .S(n5710), .Y(n4972) );
  MUX2X1 U4799 ( .B(n4976), .A(n4977), .S(n5710), .Y(n4975) );
  MUX2X1 U4800 ( .B(n4979), .A(n4980), .S(n5710), .Y(n4978) );
  MUX2X1 U4801 ( .B(n4982), .A(n4983), .S(n22), .Y(n4981) );
  MUX2X1 U4802 ( .B(n4985), .A(n4986), .S(n5710), .Y(n4984) );
  MUX2X1 U4803 ( .B(n4988), .A(n4989), .S(n5710), .Y(n4987) );
  MUX2X1 U4804 ( .B(n4991), .A(n4992), .S(n5710), .Y(n4990) );
  MUX2X1 U4805 ( .B(n4994), .A(n4995), .S(n5710), .Y(n4993) );
  MUX2X1 U4806 ( .B(n4997), .A(n4998), .S(n22), .Y(n4996) );
  MUX2X1 U4807 ( .B(n5000), .A(n5001), .S(n5711), .Y(n4999) );
  MUX2X1 U4808 ( .B(n5003), .A(n5004), .S(n5711), .Y(n5002) );
  MUX2X1 U4809 ( .B(n5006), .A(n5007), .S(n5711), .Y(n5005) );
  MUX2X1 U4810 ( .B(n5009), .A(n5010), .S(n5711), .Y(n5008) );
  MUX2X1 U4811 ( .B(n5012), .A(n5013), .S(n22), .Y(n5011) );
  MUX2X1 U4812 ( .B(n5015), .A(n5016), .S(n5711), .Y(n5014) );
  MUX2X1 U4813 ( .B(n5018), .A(n5019), .S(n5711), .Y(n5017) );
  MUX2X1 U4814 ( .B(n5021), .A(n5022), .S(n5711), .Y(n5020) );
  MUX2X1 U4815 ( .B(n5024), .A(n5025), .S(n5711), .Y(n5023) );
  MUX2X1 U4816 ( .B(n5027), .A(n5028), .S(n22), .Y(n5026) );
  MUX2X1 U4817 ( .B(n5030), .A(n5031), .S(n5711), .Y(n5029) );
  MUX2X1 U4818 ( .B(n5033), .A(n5034), .S(n5711), .Y(n5032) );
  MUX2X1 U4819 ( .B(n5036), .A(n5037), .S(n5711), .Y(n5035) );
  MUX2X1 U4820 ( .B(n5039), .A(n5040), .S(n5711), .Y(n5038) );
  MUX2X1 U4821 ( .B(n5042), .A(n5043), .S(n22), .Y(n5041) );
  MUX2X1 U4822 ( .B(n5045), .A(n5046), .S(n5712), .Y(n5044) );
  MUX2X1 U4823 ( .B(n5048), .A(n5049), .S(n5712), .Y(n5047) );
  MUX2X1 U4824 ( .B(n5051), .A(n5052), .S(n5712), .Y(n5050) );
  MUX2X1 U4825 ( .B(n5054), .A(n5055), .S(n5712), .Y(n5053) );
  MUX2X1 U4826 ( .B(n5057), .A(n5058), .S(n22), .Y(n5056) );
  MUX2X1 U4827 ( .B(n5060), .A(n5061), .S(n5712), .Y(n5059) );
  MUX2X1 U4828 ( .B(n5063), .A(n5064), .S(n5712), .Y(n5062) );
  MUX2X1 U4829 ( .B(n5066), .A(n5067), .S(n5712), .Y(n5065) );
  MUX2X1 U4830 ( .B(n5069), .A(n5070), .S(n5712), .Y(n5068) );
  MUX2X1 U4831 ( .B(n5072), .A(n5073), .S(n22), .Y(n5071) );
  MUX2X1 U4832 ( .B(n5075), .A(n5076), .S(n5712), .Y(n5074) );
  MUX2X1 U4833 ( .B(n5078), .A(n5079), .S(n5712), .Y(n5077) );
  MUX2X1 U4834 ( .B(n5081), .A(n5082), .S(n5712), .Y(n5080) );
  MUX2X1 U4835 ( .B(n5084), .A(n5085), .S(n5712), .Y(n5083) );
  MUX2X1 U4836 ( .B(n5087), .A(n5088), .S(n22), .Y(n5086) );
  MUX2X1 U4837 ( .B(n5090), .A(n5091), .S(n5713), .Y(n5089) );
  MUX2X1 U4838 ( .B(n5093), .A(n5094), .S(n5713), .Y(n5092) );
  MUX2X1 U4839 ( .B(n5096), .A(n5097), .S(n5713), .Y(n5095) );
  MUX2X1 U4840 ( .B(n5099), .A(n5100), .S(n5713), .Y(n5098) );
  MUX2X1 U4841 ( .B(n5102), .A(n5103), .S(n22), .Y(n5101) );
  MUX2X1 U4842 ( .B(n5105), .A(n5106), .S(n5713), .Y(n5104) );
  MUX2X1 U4843 ( .B(n5108), .A(n5109), .S(n5713), .Y(n5107) );
  MUX2X1 U4844 ( .B(n5111), .A(n5112), .S(n5713), .Y(n5110) );
  MUX2X1 U4845 ( .B(n5114), .A(n5115), .S(n5713), .Y(n5113) );
  MUX2X1 U4846 ( .B(n5117), .A(n5118), .S(n22), .Y(n5116) );
  MUX2X1 U4847 ( .B(n5120), .A(n5121), .S(n5713), .Y(n5119) );
  MUX2X1 U4848 ( .B(n5123), .A(n5124), .S(n5713), .Y(n5122) );
  MUX2X1 U4849 ( .B(n5126), .A(n5127), .S(n5713), .Y(n5125) );
  MUX2X1 U4850 ( .B(n5129), .A(n5130), .S(n5713), .Y(n5128) );
  MUX2X1 U4851 ( .B(n5132), .A(n5133), .S(n22), .Y(n5131) );
  MUX2X1 U4852 ( .B(n5135), .A(n5136), .S(n5714), .Y(n5134) );
  MUX2X1 U4853 ( .B(n5138), .A(n5139), .S(n5714), .Y(n5137) );
  MUX2X1 U4854 ( .B(n5141), .A(n5142), .S(n5714), .Y(n5140) );
  MUX2X1 U4855 ( .B(n5144), .A(n5145), .S(n5714), .Y(n5143) );
  MUX2X1 U4856 ( .B(n5147), .A(n5148), .S(n22), .Y(n5146) );
  MUX2X1 U4857 ( .B(n5150), .A(n5151), .S(n5714), .Y(n5149) );
  MUX2X1 U4858 ( .B(n5153), .A(n5154), .S(n5714), .Y(n5152) );
  MUX2X1 U4859 ( .B(n5156), .A(n5157), .S(n5714), .Y(n5155) );
  MUX2X1 U4860 ( .B(n5159), .A(n5160), .S(n5714), .Y(n5158) );
  MUX2X1 U4861 ( .B(n5162), .A(n5163), .S(n22), .Y(n5161) );
  MUX2X1 U4862 ( .B(n5165), .A(n5166), .S(n5714), .Y(n5164) );
  MUX2X1 U4863 ( .B(n5168), .A(n5169), .S(n5714), .Y(n5167) );
  MUX2X1 U4864 ( .B(n5171), .A(n5172), .S(n5714), .Y(n5170) );
  MUX2X1 U4865 ( .B(n5174), .A(n5175), .S(n5714), .Y(n5173) );
  MUX2X1 U4866 ( .B(n5177), .A(n5178), .S(n22), .Y(n5176) );
  MUX2X1 U4867 ( .B(n5180), .A(n5181), .S(n5715), .Y(n5179) );
  MUX2X1 U4868 ( .B(n5183), .A(n5184), .S(n5715), .Y(n5182) );
  MUX2X1 U4869 ( .B(n5186), .A(n5187), .S(n5715), .Y(n5185) );
  MUX2X1 U4870 ( .B(n5189), .A(n5190), .S(n5715), .Y(n5188) );
  MUX2X1 U4871 ( .B(n5192), .A(n5193), .S(n22), .Y(n5191) );
  MUX2X1 U4872 ( .B(n5195), .A(n5196), .S(n5715), .Y(n5194) );
  MUX2X1 U4873 ( .B(n5198), .A(n5199), .S(n5715), .Y(n5197) );
  MUX2X1 U4874 ( .B(n5201), .A(n5202), .S(n5715), .Y(n5200) );
  MUX2X1 U4875 ( .B(n5204), .A(n5205), .S(n5715), .Y(n5203) );
  MUX2X1 U4876 ( .B(n5207), .A(n5208), .S(n22), .Y(n5206) );
  MUX2X1 U4877 ( .B(n5210), .A(n5211), .S(n5715), .Y(n5209) );
  MUX2X1 U4878 ( .B(n5213), .A(n5214), .S(n5715), .Y(n5212) );
  MUX2X1 U4879 ( .B(n5216), .A(n5217), .S(n5715), .Y(n5215) );
  MUX2X1 U4880 ( .B(n5219), .A(n5220), .S(n5715), .Y(n5218) );
  MUX2X1 U4881 ( .B(n5222), .A(n5223), .S(n22), .Y(n5221) );
  MUX2X1 U4882 ( .B(n5225), .A(n5226), .S(n5716), .Y(n5224) );
  MUX2X1 U4883 ( .B(n5228), .A(n5229), .S(n5716), .Y(n5227) );
  MUX2X1 U4884 ( .B(n5231), .A(n5232), .S(n5716), .Y(n5230) );
  MUX2X1 U4885 ( .B(n5234), .A(n5235), .S(n5716), .Y(n5233) );
  MUX2X1 U4886 ( .B(n5237), .A(n5238), .S(n22), .Y(n5236) );
  MUX2X1 U4887 ( .B(n5240), .A(n5241), .S(n5716), .Y(n5239) );
  MUX2X1 U4888 ( .B(n5243), .A(n5244), .S(n5716), .Y(n5242) );
  MUX2X1 U4889 ( .B(n5246), .A(n5247), .S(n5716), .Y(n5245) );
  MUX2X1 U4890 ( .B(n5249), .A(n5250), .S(n5716), .Y(n5248) );
  MUX2X1 U4891 ( .B(n5252), .A(n5253), .S(n22), .Y(n5251) );
  MUX2X1 U4892 ( .B(n5255), .A(n5256), .S(n5716), .Y(n5254) );
  MUX2X1 U4893 ( .B(n5258), .A(n5259), .S(n5716), .Y(n5257) );
  MUX2X1 U4894 ( .B(n5261), .A(n5262), .S(n5716), .Y(n5260) );
  MUX2X1 U4895 ( .B(n5264), .A(n5265), .S(n5716), .Y(n5263) );
  MUX2X1 U4896 ( .B(n5267), .A(n5268), .S(n22), .Y(n5266) );
  MUX2X1 U4897 ( .B(n5270), .A(n5271), .S(n5717), .Y(n5269) );
  MUX2X1 U4898 ( .B(n5273), .A(n5274), .S(n5717), .Y(n5272) );
  MUX2X1 U4899 ( .B(n5276), .A(n5277), .S(n5717), .Y(n5275) );
  MUX2X1 U4900 ( .B(n5279), .A(n5280), .S(n5717), .Y(n5278) );
  MUX2X1 U4901 ( .B(n5282), .A(n5283), .S(n22), .Y(n5281) );
  MUX2X1 U4902 ( .B(n5285), .A(n5286), .S(n5717), .Y(n5284) );
  MUX2X1 U4903 ( .B(n5288), .A(n5289), .S(n5717), .Y(n5287) );
  MUX2X1 U4904 ( .B(n5291), .A(n5292), .S(n5717), .Y(n5290) );
  MUX2X1 U4905 ( .B(n5294), .A(n5295), .S(n5717), .Y(n5293) );
  MUX2X1 U4906 ( .B(n5297), .A(n5298), .S(n22), .Y(n5296) );
  MUX2X1 U4907 ( .B(n5300), .A(n5301), .S(n5717), .Y(n5299) );
  MUX2X1 U4908 ( .B(n5303), .A(n5304), .S(n5717), .Y(n5302) );
  MUX2X1 U4909 ( .B(n5306), .A(n5307), .S(n5717), .Y(n5305) );
  MUX2X1 U4910 ( .B(n5309), .A(n5310), .S(n5717), .Y(n5308) );
  MUX2X1 U4911 ( .B(n5312), .A(n5313), .S(n22), .Y(n5311) );
  MUX2X1 U4912 ( .B(n5315), .A(n5316), .S(n5718), .Y(n5314) );
  MUX2X1 U4913 ( .B(n5318), .A(n5319), .S(n5718), .Y(n5317) );
  MUX2X1 U4914 ( .B(n5321), .A(n5322), .S(n5718), .Y(n5320) );
  MUX2X1 U4915 ( .B(n5324), .A(n5325), .S(n5718), .Y(n5323) );
  MUX2X1 U4916 ( .B(n5327), .A(n5328), .S(n22), .Y(n5326) );
  MUX2X1 U4917 ( .B(n5330), .A(n5331), .S(n5718), .Y(n5329) );
  MUX2X1 U4918 ( .B(n5333), .A(n5334), .S(n5718), .Y(n5332) );
  MUX2X1 U4919 ( .B(n5336), .A(n5337), .S(n5718), .Y(n5335) );
  MUX2X1 U4920 ( .B(n5339), .A(n5340), .S(n5718), .Y(n5338) );
  MUX2X1 U4921 ( .B(n5342), .A(n5343), .S(n22), .Y(n5341) );
  MUX2X1 U4922 ( .B(n5345), .A(n5346), .S(n5718), .Y(n5344) );
  MUX2X1 U4923 ( .B(n5348), .A(n5349), .S(n5718), .Y(n5347) );
  MUX2X1 U4924 ( .B(n5351), .A(n5352), .S(n5718), .Y(n5350) );
  MUX2X1 U4925 ( .B(n5354), .A(n5355), .S(n5718), .Y(n5353) );
  MUX2X1 U4926 ( .B(n5357), .A(n5358), .S(n22), .Y(n5356) );
  MUX2X1 U4927 ( .B(n5360), .A(n5361), .S(n5719), .Y(n5359) );
  MUX2X1 U4928 ( .B(n5363), .A(n5364), .S(n5719), .Y(n5362) );
  MUX2X1 U4929 ( .B(n5366), .A(n5367), .S(n5719), .Y(n5365) );
  MUX2X1 U4930 ( .B(n5369), .A(n5370), .S(n5719), .Y(n5368) );
  MUX2X1 U4931 ( .B(n5372), .A(n5373), .S(n22), .Y(n5371) );
  MUX2X1 U4932 ( .B(n5375), .A(n5376), .S(n5719), .Y(n5374) );
  MUX2X1 U4933 ( .B(n5378), .A(n5379), .S(n5719), .Y(n5377) );
  MUX2X1 U4934 ( .B(n5381), .A(n5382), .S(n5719), .Y(n5380) );
  MUX2X1 U4935 ( .B(n5384), .A(n5385), .S(n5719), .Y(n5383) );
  MUX2X1 U4936 ( .B(n5387), .A(n5388), .S(n22), .Y(n5386) );
  MUX2X1 U4937 ( .B(n5390), .A(n5391), .S(n5719), .Y(n5389) );
  MUX2X1 U4938 ( .B(n5393), .A(n5394), .S(n5719), .Y(n5392) );
  MUX2X1 U4939 ( .B(n5396), .A(n5397), .S(n5719), .Y(n5395) );
  MUX2X1 U4940 ( .B(n5399), .A(n5400), .S(n5719), .Y(n5398) );
  MUX2X1 U4941 ( .B(n5402), .A(n5403), .S(n22), .Y(n5401) );
  MUX2X1 U4942 ( .B(n5405), .A(n5406), .S(n5720), .Y(n5404) );
  MUX2X1 U4943 ( .B(n5408), .A(n5409), .S(n5720), .Y(n5407) );
  MUX2X1 U4944 ( .B(n5411), .A(n5412), .S(n5720), .Y(n5410) );
  MUX2X1 U4945 ( .B(n5414), .A(n5415), .S(n5720), .Y(n5413) );
  MUX2X1 U4946 ( .B(n5417), .A(n5418), .S(n22), .Y(n5416) );
  MUX2X1 U4947 ( .B(n5420), .A(n5421), .S(n5720), .Y(n5419) );
  MUX2X1 U4948 ( .B(n5423), .A(n5424), .S(n5720), .Y(n5422) );
  MUX2X1 U4949 ( .B(n5426), .A(n5427), .S(n5720), .Y(n5425) );
  MUX2X1 U4950 ( .B(n5429), .A(n5430), .S(n5720), .Y(n5428) );
  MUX2X1 U4951 ( .B(n5432), .A(n5433), .S(n22), .Y(n5431) );
  MUX2X1 U4952 ( .B(n5435), .A(n5436), .S(n5720), .Y(n5434) );
  MUX2X1 U4953 ( .B(n5438), .A(n5439), .S(n5720), .Y(n5437) );
  MUX2X1 U4954 ( .B(n5441), .A(n5442), .S(n5720), .Y(n5440) );
  MUX2X1 U4955 ( .B(n5444), .A(n5445), .S(n5720), .Y(n5443) );
  MUX2X1 U4956 ( .B(n5447), .A(n5448), .S(n22), .Y(n5446) );
  MUX2X1 U4957 ( .B(n5450), .A(n5451), .S(n5721), .Y(n5449) );
  MUX2X1 U4958 ( .B(n5453), .A(n5454), .S(n5721), .Y(n5452) );
  MUX2X1 U4959 ( .B(n5456), .A(n5457), .S(n5721), .Y(n5455) );
  MUX2X1 U4960 ( .B(n5459), .A(n5460), .S(n5721), .Y(n5458) );
  MUX2X1 U4961 ( .B(n5462), .A(n5463), .S(n22), .Y(n5461) );
  MUX2X1 U4962 ( .B(n5465), .A(n5466), .S(n5721), .Y(n5464) );
  MUX2X1 U4963 ( .B(n5468), .A(n5469), .S(n5721), .Y(n5467) );
  MUX2X1 U4964 ( .B(n5471), .A(n5472), .S(n5721), .Y(n5470) );
  MUX2X1 U4965 ( .B(n5474), .A(n5475), .S(n5721), .Y(n5473) );
  MUX2X1 U4966 ( .B(n5477), .A(n5478), .S(n22), .Y(n5476) );
  MUX2X1 U4967 ( .B(n5480), .A(n5481), .S(n5721), .Y(n5479) );
  MUX2X1 U4968 ( .B(n5483), .A(n5484), .S(n5721), .Y(n5482) );
  MUX2X1 U4969 ( .B(n5486), .A(n5487), .S(n5721), .Y(n5485) );
  MUX2X1 U4970 ( .B(n5489), .A(n5490), .S(n5721), .Y(n5488) );
  MUX2X1 U4971 ( .B(n5492), .A(n5493), .S(n22), .Y(n5491) );
  MUX2X1 U4972 ( .B(n5495), .A(n5496), .S(n5722), .Y(n5494) );
  MUX2X1 U4973 ( .B(n5498), .A(n5499), .S(n5722), .Y(n5497) );
  MUX2X1 U4974 ( .B(n5501), .A(n5502), .S(n5722), .Y(n5500) );
  MUX2X1 U4975 ( .B(n5504), .A(n5505), .S(n5722), .Y(n5503) );
  MUX2X1 U4976 ( .B(n5507), .A(n5508), .S(n22), .Y(n5506) );
  MUX2X1 U4977 ( .B(n5510), .A(n5511), .S(n5722), .Y(n5509) );
  MUX2X1 U4978 ( .B(n5513), .A(n5514), .S(n5722), .Y(n5512) );
  MUX2X1 U4979 ( .B(n5516), .A(n5517), .S(n5722), .Y(n5515) );
  MUX2X1 U4980 ( .B(n5519), .A(n5520), .S(n5722), .Y(n5518) );
  MUX2X1 U4981 ( .B(n5522), .A(n5523), .S(n22), .Y(n5521) );
  MUX2X1 U4982 ( .B(n5525), .A(n5526), .S(n5722), .Y(n5524) );
  MUX2X1 U4983 ( .B(n5528), .A(n5529), .S(n5722), .Y(n5527) );
  MUX2X1 U4984 ( .B(n5531), .A(n5532), .S(n5722), .Y(n5530) );
  MUX2X1 U4985 ( .B(n5534), .A(n5535), .S(n5722), .Y(n5533) );
  MUX2X1 U4986 ( .B(n5537), .A(n5538), .S(n22), .Y(n5536) );
  MUX2X1 U4987 ( .B(n5540), .A(n5541), .S(n5723), .Y(n5539) );
  MUX2X1 U4988 ( .B(n5543), .A(n5544), .S(n5723), .Y(n5542) );
  MUX2X1 U4989 ( .B(n5546), .A(n5547), .S(n5723), .Y(n5545) );
  MUX2X1 U4990 ( .B(n5549), .A(n5550), .S(n5723), .Y(n5548) );
  MUX2X1 U4991 ( .B(n5552), .A(n5553), .S(n22), .Y(n5551) );
  MUX2X1 U4992 ( .B(n5555), .A(n5556), .S(n5723), .Y(n5554) );
  MUX2X1 U4993 ( .B(n5558), .A(n5559), .S(n5723), .Y(n5557) );
  MUX2X1 U4994 ( .B(n5561), .A(n5562), .S(n5723), .Y(n5560) );
  MUX2X1 U4995 ( .B(n5564), .A(n5565), .S(n5723), .Y(n5563) );
  MUX2X1 U4996 ( .B(n5567), .A(n5568), .S(n22), .Y(n5566) );
  MUX2X1 U4997 ( .B(n5570), .A(n5571), .S(n5723), .Y(n5569) );
  MUX2X1 U4998 ( .B(n5573), .A(n5574), .S(n5723), .Y(n5572) );
  MUX2X1 U4999 ( .B(n5576), .A(n5577), .S(n5723), .Y(n5575) );
  MUX2X1 U5000 ( .B(n5579), .A(n5580), .S(n5723), .Y(n5578) );
  MUX2X1 U5001 ( .B(n5582), .A(n5583), .S(n22), .Y(n5581) );
  MUX2X1 U5002 ( .B(fifo_array[1260]), .A(fifo_array[1302]), .S(n5638), .Y(
        n4326) );
  MUX2X1 U5003 ( .B(fifo_array[1176]), .A(fifo_array[1218]), .S(n5638), .Y(
        n4325) );
  MUX2X1 U5004 ( .B(fifo_array[1092]), .A(fifo_array[1134]), .S(n5638), .Y(
        n4329) );
  MUX2X1 U5005 ( .B(fifo_array[1008]), .A(fifo_array[1050]), .S(n5638), .Y(
        n4328) );
  MUX2X1 U5006 ( .B(n4327), .A(n4324), .S(n5724), .Y(n4338) );
  MUX2X1 U5007 ( .B(fifo_array[924]), .A(fifo_array[966]), .S(n5638), .Y(n4332) );
  MUX2X1 U5008 ( .B(fifo_array[840]), .A(fifo_array[882]), .S(n5638), .Y(n4331) );
  MUX2X1 U5009 ( .B(fifo_array[756]), .A(fifo_array[798]), .S(n5638), .Y(n4335) );
  MUX2X1 U5010 ( .B(fifo_array[672]), .A(fifo_array[714]), .S(n5638), .Y(n4334) );
  MUX2X1 U5011 ( .B(n4333), .A(n4330), .S(n5724), .Y(n4337) );
  MUX2X1 U5012 ( .B(fifo_array[588]), .A(fifo_array[630]), .S(n5638), .Y(n4341) );
  MUX2X1 U5013 ( .B(fifo_array[504]), .A(fifo_array[546]), .S(n5638), .Y(n4340) );
  MUX2X1 U5014 ( .B(fifo_array[420]), .A(fifo_array[462]), .S(n5638), .Y(n4344) );
  MUX2X1 U5015 ( .B(fifo_array[336]), .A(fifo_array[378]), .S(n5638), .Y(n4343) );
  MUX2X1 U5016 ( .B(n4342), .A(n4339), .S(n5724), .Y(n4353) );
  MUX2X1 U5017 ( .B(fifo_array[252]), .A(fifo_array[294]), .S(n5639), .Y(n4347) );
  MUX2X1 U5018 ( .B(fifo_array[168]), .A(fifo_array[210]), .S(n5639), .Y(n4346) );
  MUX2X1 U5019 ( .B(fifo_array[84]), .A(fifo_array[126]), .S(n5639), .Y(n4350)
         );
  MUX2X1 U5020 ( .B(fifo_array[0]), .A(fifo_array[42]), .S(n5639), .Y(n4349)
         );
  MUX2X1 U5021 ( .B(n4348), .A(n4345), .S(n5724), .Y(n4352) );
  MUX2X1 U5022 ( .B(n4351), .A(n4336), .S(n23), .Y(n5584) );
  MUX2X1 U5023 ( .B(fifo_array[1261]), .A(fifo_array[1303]), .S(n5639), .Y(
        n4356) );
  MUX2X1 U5024 ( .B(fifo_array[1177]), .A(fifo_array[1219]), .S(n5639), .Y(
        n4355) );
  MUX2X1 U5025 ( .B(fifo_array[1093]), .A(fifo_array[1135]), .S(n5639), .Y(
        n4359) );
  MUX2X1 U5026 ( .B(fifo_array[1009]), .A(fifo_array[1051]), .S(n5639), .Y(
        n4358) );
  MUX2X1 U5027 ( .B(n4357), .A(n4354), .S(n5724), .Y(n4368) );
  MUX2X1 U5028 ( .B(fifo_array[925]), .A(fifo_array[967]), .S(n5639), .Y(n4362) );
  MUX2X1 U5029 ( .B(fifo_array[841]), .A(fifo_array[883]), .S(n5639), .Y(n4361) );
  MUX2X1 U5030 ( .B(fifo_array[757]), .A(fifo_array[799]), .S(n5639), .Y(n4365) );
  MUX2X1 U5031 ( .B(fifo_array[673]), .A(fifo_array[715]), .S(n5639), .Y(n4364) );
  MUX2X1 U5032 ( .B(n4363), .A(n4360), .S(n5724), .Y(n4367) );
  MUX2X1 U5033 ( .B(fifo_array[589]), .A(fifo_array[631]), .S(n5640), .Y(n4371) );
  MUX2X1 U5034 ( .B(fifo_array[505]), .A(fifo_array[547]), .S(n5640), .Y(n4370) );
  MUX2X1 U5035 ( .B(fifo_array[421]), .A(fifo_array[463]), .S(n5640), .Y(n4374) );
  MUX2X1 U5036 ( .B(fifo_array[337]), .A(fifo_array[379]), .S(n5640), .Y(n4373) );
  MUX2X1 U5037 ( .B(n4372), .A(n4369), .S(n5724), .Y(n4383) );
  MUX2X1 U5038 ( .B(fifo_array[253]), .A(fifo_array[295]), .S(n5640), .Y(n4377) );
  MUX2X1 U5039 ( .B(fifo_array[169]), .A(fifo_array[211]), .S(n5640), .Y(n4376) );
  MUX2X1 U5040 ( .B(fifo_array[85]), .A(fifo_array[127]), .S(n5640), .Y(n4380)
         );
  MUX2X1 U5041 ( .B(fifo_array[1]), .A(fifo_array[43]), .S(n5640), .Y(n4379)
         );
  MUX2X1 U5042 ( .B(n4378), .A(n4375), .S(n5724), .Y(n4382) );
  MUX2X1 U5043 ( .B(n4381), .A(n4366), .S(n23), .Y(n5585) );
  MUX2X1 U5044 ( .B(fifo_array[1262]), .A(fifo_array[1304]), .S(n5640), .Y(
        n4386) );
  MUX2X1 U5045 ( .B(fifo_array[1178]), .A(fifo_array[1220]), .S(n5640), .Y(
        n4385) );
  MUX2X1 U5046 ( .B(fifo_array[1094]), .A(fifo_array[1136]), .S(n5640), .Y(
        n4389) );
  MUX2X1 U5047 ( .B(fifo_array[1010]), .A(fifo_array[1052]), .S(n5640), .Y(
        n4388) );
  MUX2X1 U5048 ( .B(n4387), .A(n4384), .S(n5724), .Y(n4398) );
  MUX2X1 U5049 ( .B(fifo_array[926]), .A(fifo_array[968]), .S(n5641), .Y(n4392) );
  MUX2X1 U5050 ( .B(fifo_array[842]), .A(fifo_array[884]), .S(n5641), .Y(n4391) );
  MUX2X1 U5051 ( .B(fifo_array[758]), .A(fifo_array[800]), .S(n5641), .Y(n4395) );
  MUX2X1 U5052 ( .B(fifo_array[674]), .A(fifo_array[716]), .S(n5641), .Y(n4394) );
  MUX2X1 U5053 ( .B(n4393), .A(n4390), .S(n5724), .Y(n4397) );
  MUX2X1 U5054 ( .B(fifo_array[590]), .A(fifo_array[632]), .S(n5641), .Y(n4401) );
  MUX2X1 U5055 ( .B(fifo_array[506]), .A(fifo_array[548]), .S(n5641), .Y(n4400) );
  MUX2X1 U5056 ( .B(fifo_array[422]), .A(fifo_array[464]), .S(n5641), .Y(n4404) );
  MUX2X1 U5057 ( .B(fifo_array[338]), .A(fifo_array[380]), .S(n5641), .Y(n4403) );
  MUX2X1 U5058 ( .B(n4402), .A(n4399), .S(n5724), .Y(n4413) );
  MUX2X1 U5059 ( .B(fifo_array[254]), .A(fifo_array[296]), .S(n5641), .Y(n4407) );
  MUX2X1 U5060 ( .B(fifo_array[170]), .A(fifo_array[212]), .S(n5641), .Y(n4406) );
  MUX2X1 U5061 ( .B(fifo_array[86]), .A(fifo_array[128]), .S(n5641), .Y(n4410)
         );
  MUX2X1 U5062 ( .B(fifo_array[2]), .A(fifo_array[44]), .S(n5641), .Y(n4409)
         );
  MUX2X1 U5063 ( .B(n4408), .A(n4405), .S(n5724), .Y(n4412) );
  MUX2X1 U5064 ( .B(n4411), .A(n4396), .S(n23), .Y(n5586) );
  MUX2X1 U5065 ( .B(fifo_array[1263]), .A(fifo_array[1305]), .S(n5642), .Y(
        n4416) );
  MUX2X1 U5066 ( .B(fifo_array[1179]), .A(fifo_array[1221]), .S(n5642), .Y(
        n4415) );
  MUX2X1 U5067 ( .B(fifo_array[1095]), .A(fifo_array[1137]), .S(n5642), .Y(
        n4419) );
  MUX2X1 U5068 ( .B(fifo_array[1011]), .A(fifo_array[1053]), .S(n5642), .Y(
        n4418) );
  MUX2X1 U5069 ( .B(n4417), .A(n4414), .S(n5725), .Y(n4428) );
  MUX2X1 U5070 ( .B(fifo_array[927]), .A(fifo_array[969]), .S(n5642), .Y(n4422) );
  MUX2X1 U5071 ( .B(fifo_array[843]), .A(fifo_array[885]), .S(n5642), .Y(n4421) );
  MUX2X1 U5072 ( .B(fifo_array[759]), .A(fifo_array[801]), .S(n5642), .Y(n4425) );
  MUX2X1 U5073 ( .B(fifo_array[675]), .A(fifo_array[717]), .S(n5642), .Y(n4424) );
  MUX2X1 U5074 ( .B(n4423), .A(n4420), .S(n5725), .Y(n4427) );
  MUX2X1 U5075 ( .B(fifo_array[591]), .A(fifo_array[633]), .S(n5642), .Y(n4431) );
  MUX2X1 U5076 ( .B(fifo_array[507]), .A(fifo_array[549]), .S(n5642), .Y(n4430) );
  MUX2X1 U5077 ( .B(fifo_array[423]), .A(fifo_array[465]), .S(n5642), .Y(n4434) );
  MUX2X1 U5078 ( .B(fifo_array[339]), .A(fifo_array[381]), .S(n5642), .Y(n4433) );
  MUX2X1 U5079 ( .B(n4432), .A(n4429), .S(n5725), .Y(n4443) );
  MUX2X1 U5080 ( .B(fifo_array[255]), .A(fifo_array[297]), .S(n5643), .Y(n4437) );
  MUX2X1 U5081 ( .B(fifo_array[171]), .A(fifo_array[213]), .S(n5643), .Y(n4436) );
  MUX2X1 U5082 ( .B(fifo_array[87]), .A(fifo_array[129]), .S(n5643), .Y(n4440)
         );
  MUX2X1 U5083 ( .B(fifo_array[3]), .A(fifo_array[45]), .S(n5643), .Y(n4439)
         );
  MUX2X1 U5084 ( .B(n4438), .A(n4435), .S(n5725), .Y(n4442) );
  MUX2X1 U5085 ( .B(n4441), .A(n4426), .S(n23), .Y(n5587) );
  MUX2X1 U5086 ( .B(fifo_array[1264]), .A(fifo_array[1306]), .S(n5643), .Y(
        n4446) );
  MUX2X1 U5087 ( .B(fifo_array[1180]), .A(fifo_array[1222]), .S(n5643), .Y(
        n4445) );
  MUX2X1 U5088 ( .B(fifo_array[1096]), .A(fifo_array[1138]), .S(n5643), .Y(
        n4449) );
  MUX2X1 U5089 ( .B(fifo_array[1012]), .A(fifo_array[1054]), .S(n5643), .Y(
        n4448) );
  MUX2X1 U5090 ( .B(n4447), .A(n4444), .S(n5725), .Y(n4458) );
  MUX2X1 U5091 ( .B(fifo_array[928]), .A(fifo_array[970]), .S(n5643), .Y(n4452) );
  MUX2X1 U5092 ( .B(fifo_array[844]), .A(fifo_array[886]), .S(n5643), .Y(n4451) );
  MUX2X1 U5093 ( .B(fifo_array[760]), .A(fifo_array[802]), .S(n5643), .Y(n4455) );
  MUX2X1 U5094 ( .B(fifo_array[676]), .A(fifo_array[718]), .S(n5643), .Y(n4454) );
  MUX2X1 U5095 ( .B(n4453), .A(n4450), .S(n5725), .Y(n4457) );
  MUX2X1 U5096 ( .B(fifo_array[592]), .A(fifo_array[634]), .S(n5644), .Y(n4461) );
  MUX2X1 U5097 ( .B(fifo_array[508]), .A(fifo_array[550]), .S(n5644), .Y(n4460) );
  MUX2X1 U5098 ( .B(fifo_array[424]), .A(fifo_array[466]), .S(n5644), .Y(n4464) );
  MUX2X1 U5099 ( .B(fifo_array[340]), .A(fifo_array[382]), .S(n5644), .Y(n4463) );
  MUX2X1 U5100 ( .B(n4462), .A(n4459), .S(n5725), .Y(n4473) );
  MUX2X1 U5101 ( .B(fifo_array[256]), .A(fifo_array[298]), .S(n5644), .Y(n4467) );
  MUX2X1 U5102 ( .B(fifo_array[172]), .A(fifo_array[214]), .S(n5644), .Y(n4466) );
  MUX2X1 U5103 ( .B(fifo_array[88]), .A(fifo_array[130]), .S(n5644), .Y(n4470)
         );
  MUX2X1 U5104 ( .B(fifo_array[4]), .A(fifo_array[46]), .S(n5644), .Y(n4469)
         );
  MUX2X1 U5105 ( .B(n4468), .A(n4465), .S(n5725), .Y(n4472) );
  MUX2X1 U5106 ( .B(n4471), .A(n4456), .S(n23), .Y(n5588) );
  MUX2X1 U5107 ( .B(fifo_array[1265]), .A(fifo_array[1307]), .S(n5644), .Y(
        n4476) );
  MUX2X1 U5108 ( .B(fifo_array[1181]), .A(fifo_array[1223]), .S(n5644), .Y(
        n4475) );
  MUX2X1 U5109 ( .B(fifo_array[1097]), .A(fifo_array[1139]), .S(n5644), .Y(
        n4479) );
  MUX2X1 U5110 ( .B(fifo_array[1013]), .A(fifo_array[1055]), .S(n5644), .Y(
        n4478) );
  MUX2X1 U5111 ( .B(n4477), .A(n4474), .S(n5725), .Y(n4488) );
  MUX2X1 U5112 ( .B(fifo_array[929]), .A(fifo_array[971]), .S(n5645), .Y(n4482) );
  MUX2X1 U5113 ( .B(fifo_array[845]), .A(fifo_array[887]), .S(n5645), .Y(n4481) );
  MUX2X1 U5114 ( .B(fifo_array[761]), .A(fifo_array[803]), .S(n5645), .Y(n4485) );
  MUX2X1 U5115 ( .B(fifo_array[677]), .A(fifo_array[719]), .S(n5645), .Y(n4484) );
  MUX2X1 U5116 ( .B(n4483), .A(n4480), .S(n5725), .Y(n4487) );
  MUX2X1 U5117 ( .B(fifo_array[593]), .A(fifo_array[635]), .S(n5645), .Y(n4491) );
  MUX2X1 U5118 ( .B(fifo_array[509]), .A(fifo_array[551]), .S(n5645), .Y(n4490) );
  MUX2X1 U5119 ( .B(fifo_array[425]), .A(fifo_array[467]), .S(n5645), .Y(n4494) );
  MUX2X1 U5120 ( .B(fifo_array[341]), .A(fifo_array[383]), .S(n5645), .Y(n4493) );
  MUX2X1 U5121 ( .B(n4492), .A(n4489), .S(n5725), .Y(n4503) );
  MUX2X1 U5122 ( .B(fifo_array[257]), .A(fifo_array[299]), .S(n5645), .Y(n4497) );
  MUX2X1 U5123 ( .B(fifo_array[173]), .A(fifo_array[215]), .S(n5645), .Y(n4496) );
  MUX2X1 U5124 ( .B(fifo_array[89]), .A(fifo_array[131]), .S(n5645), .Y(n4500)
         );
  MUX2X1 U5125 ( .B(fifo_array[5]), .A(fifo_array[47]), .S(n5645), .Y(n4499)
         );
  MUX2X1 U5126 ( .B(n4498), .A(n4495), .S(n5725), .Y(n4502) );
  MUX2X1 U5127 ( .B(n4501), .A(n4486), .S(n23), .Y(n5589) );
  MUX2X1 U5128 ( .B(fifo_array[1266]), .A(fifo_array[1308]), .S(n5646), .Y(
        n4506) );
  MUX2X1 U5129 ( .B(fifo_array[1182]), .A(fifo_array[1224]), .S(n5646), .Y(
        n4505) );
  MUX2X1 U5130 ( .B(fifo_array[1098]), .A(fifo_array[1140]), .S(n5646), .Y(
        n4509) );
  MUX2X1 U5131 ( .B(fifo_array[1014]), .A(fifo_array[1056]), .S(n5646), .Y(
        n4508) );
  MUX2X1 U5132 ( .B(n4507), .A(n4504), .S(n5726), .Y(n4518) );
  MUX2X1 U5133 ( .B(fifo_array[930]), .A(fifo_array[972]), .S(n5646), .Y(n4512) );
  MUX2X1 U5134 ( .B(fifo_array[846]), .A(fifo_array[888]), .S(n5646), .Y(n4511) );
  MUX2X1 U5135 ( .B(fifo_array[762]), .A(fifo_array[804]), .S(n5646), .Y(n4515) );
  MUX2X1 U5136 ( .B(fifo_array[678]), .A(fifo_array[720]), .S(n5646), .Y(n4514) );
  MUX2X1 U5137 ( .B(n4513), .A(n4510), .S(n5726), .Y(n4517) );
  MUX2X1 U5138 ( .B(fifo_array[594]), .A(fifo_array[636]), .S(n5646), .Y(n4521) );
  MUX2X1 U5139 ( .B(fifo_array[510]), .A(fifo_array[552]), .S(n5646), .Y(n4520) );
  MUX2X1 U5140 ( .B(fifo_array[426]), .A(fifo_array[468]), .S(n5646), .Y(n4524) );
  MUX2X1 U5141 ( .B(fifo_array[342]), .A(fifo_array[384]), .S(n5646), .Y(n4523) );
  MUX2X1 U5142 ( .B(n4522), .A(n4519), .S(n5726), .Y(n4533) );
  MUX2X1 U5143 ( .B(fifo_array[258]), .A(fifo_array[300]), .S(n5647), .Y(n4527) );
  MUX2X1 U5144 ( .B(fifo_array[174]), .A(fifo_array[216]), .S(n5647), .Y(n4526) );
  MUX2X1 U5145 ( .B(fifo_array[90]), .A(fifo_array[132]), .S(n5647), .Y(n4530)
         );
  MUX2X1 U5146 ( .B(fifo_array[6]), .A(fifo_array[48]), .S(n5647), .Y(n4529)
         );
  MUX2X1 U5147 ( .B(n4528), .A(n4525), .S(n5726), .Y(n4532) );
  MUX2X1 U5148 ( .B(n4531), .A(n4516), .S(n23), .Y(n5590) );
  MUX2X1 U5149 ( .B(fifo_array[1267]), .A(fifo_array[1309]), .S(n5647), .Y(
        n4536) );
  MUX2X1 U5150 ( .B(fifo_array[1183]), .A(fifo_array[1225]), .S(n5647), .Y(
        n4535) );
  MUX2X1 U5151 ( .B(fifo_array[1099]), .A(fifo_array[1141]), .S(n5647), .Y(
        n4539) );
  MUX2X1 U5152 ( .B(fifo_array[1015]), .A(fifo_array[1057]), .S(n5647), .Y(
        n4538) );
  MUX2X1 U5153 ( .B(n4537), .A(n4534), .S(n5726), .Y(n4548) );
  MUX2X1 U5154 ( .B(fifo_array[931]), .A(fifo_array[973]), .S(n5647), .Y(n4542) );
  MUX2X1 U5155 ( .B(fifo_array[847]), .A(fifo_array[889]), .S(n5647), .Y(n4541) );
  MUX2X1 U5156 ( .B(fifo_array[763]), .A(fifo_array[805]), .S(n5647), .Y(n4545) );
  MUX2X1 U5157 ( .B(fifo_array[679]), .A(fifo_array[721]), .S(n5647), .Y(n4544) );
  MUX2X1 U5158 ( .B(n4543), .A(n4540), .S(n5726), .Y(n4547) );
  MUX2X1 U5159 ( .B(fifo_array[595]), .A(fifo_array[637]), .S(n5648), .Y(n4551) );
  MUX2X1 U5160 ( .B(fifo_array[511]), .A(fifo_array[553]), .S(n5648), .Y(n4550) );
  MUX2X1 U5161 ( .B(fifo_array[427]), .A(fifo_array[469]), .S(n5648), .Y(n4554) );
  MUX2X1 U5162 ( .B(fifo_array[343]), .A(fifo_array[385]), .S(n5648), .Y(n4553) );
  MUX2X1 U5163 ( .B(n4552), .A(n4549), .S(n5726), .Y(n4563) );
  MUX2X1 U5164 ( .B(fifo_array[259]), .A(fifo_array[301]), .S(n5648), .Y(n4557) );
  MUX2X1 U5165 ( .B(fifo_array[175]), .A(fifo_array[217]), .S(n5648), .Y(n4556) );
  MUX2X1 U5166 ( .B(fifo_array[91]), .A(fifo_array[133]), .S(n5648), .Y(n4560)
         );
  MUX2X1 U5167 ( .B(fifo_array[7]), .A(fifo_array[49]), .S(n5648), .Y(n4559)
         );
  MUX2X1 U5168 ( .B(n4558), .A(n4555), .S(n5726), .Y(n4562) );
  MUX2X1 U5169 ( .B(n4561), .A(n4546), .S(n23), .Y(n5591) );
  MUX2X1 U5170 ( .B(fifo_array[1268]), .A(fifo_array[1310]), .S(n5648), .Y(
        n4566) );
  MUX2X1 U5171 ( .B(fifo_array[1184]), .A(fifo_array[1226]), .S(n5648), .Y(
        n4565) );
  MUX2X1 U5172 ( .B(fifo_array[1100]), .A(fifo_array[1142]), .S(n5648), .Y(
        n4569) );
  MUX2X1 U5173 ( .B(fifo_array[1016]), .A(fifo_array[1058]), .S(n5648), .Y(
        n4568) );
  MUX2X1 U5174 ( .B(n4567), .A(n4564), .S(n5726), .Y(n4578) );
  MUX2X1 U5175 ( .B(fifo_array[932]), .A(fifo_array[974]), .S(n5649), .Y(n4572) );
  MUX2X1 U5176 ( .B(fifo_array[848]), .A(fifo_array[890]), .S(n5649), .Y(n4571) );
  MUX2X1 U5177 ( .B(fifo_array[764]), .A(fifo_array[806]), .S(n5649), .Y(n4575) );
  MUX2X1 U5178 ( .B(fifo_array[680]), .A(fifo_array[722]), .S(n5649), .Y(n4574) );
  MUX2X1 U5179 ( .B(n4573), .A(n4570), .S(n5726), .Y(n4577) );
  MUX2X1 U5180 ( .B(fifo_array[596]), .A(fifo_array[638]), .S(n5649), .Y(n4581) );
  MUX2X1 U5181 ( .B(fifo_array[512]), .A(fifo_array[554]), .S(n5649), .Y(n4580) );
  MUX2X1 U5182 ( .B(fifo_array[428]), .A(fifo_array[470]), .S(n5649), .Y(n4584) );
  MUX2X1 U5183 ( .B(fifo_array[344]), .A(fifo_array[386]), .S(n5649), .Y(n4583) );
  MUX2X1 U5184 ( .B(n4582), .A(n4579), .S(n5726), .Y(n4593) );
  MUX2X1 U5185 ( .B(fifo_array[260]), .A(fifo_array[302]), .S(n5649), .Y(n4587) );
  MUX2X1 U5186 ( .B(fifo_array[176]), .A(fifo_array[218]), .S(n5649), .Y(n4586) );
  MUX2X1 U5187 ( .B(fifo_array[92]), .A(fifo_array[134]), .S(n5649), .Y(n4590)
         );
  MUX2X1 U5188 ( .B(fifo_array[8]), .A(fifo_array[50]), .S(n5649), .Y(n4589)
         );
  MUX2X1 U5189 ( .B(n4588), .A(n4585), .S(n5726), .Y(n4592) );
  MUX2X1 U5190 ( .B(n4591), .A(n4576), .S(n23), .Y(n5592) );
  MUX2X1 U5191 ( .B(fifo_array[1269]), .A(fifo_array[1311]), .S(n5650), .Y(
        n4596) );
  MUX2X1 U5192 ( .B(fifo_array[1185]), .A(fifo_array[1227]), .S(n5650), .Y(
        n4595) );
  MUX2X1 U5193 ( .B(fifo_array[1101]), .A(fifo_array[1143]), .S(n5650), .Y(
        n4599) );
  MUX2X1 U5194 ( .B(fifo_array[1017]), .A(fifo_array[1059]), .S(n5650), .Y(
        n4598) );
  MUX2X1 U5195 ( .B(n4597), .A(n4594), .S(n5727), .Y(n4608) );
  MUX2X1 U5196 ( .B(fifo_array[933]), .A(fifo_array[975]), .S(n5650), .Y(n4602) );
  MUX2X1 U5197 ( .B(fifo_array[849]), .A(fifo_array[891]), .S(n5650), .Y(n4601) );
  MUX2X1 U5198 ( .B(fifo_array[765]), .A(fifo_array[807]), .S(n5650), .Y(n4605) );
  MUX2X1 U5199 ( .B(fifo_array[681]), .A(fifo_array[723]), .S(n5650), .Y(n4604) );
  MUX2X1 U5200 ( .B(n4603), .A(n4600), .S(n5727), .Y(n4607) );
  MUX2X1 U5201 ( .B(fifo_array[597]), .A(fifo_array[639]), .S(n5650), .Y(n4611) );
  MUX2X1 U5202 ( .B(fifo_array[513]), .A(fifo_array[555]), .S(n5650), .Y(n4610) );
  MUX2X1 U5203 ( .B(fifo_array[429]), .A(fifo_array[471]), .S(n5650), .Y(n4614) );
  MUX2X1 U5204 ( .B(fifo_array[345]), .A(fifo_array[387]), .S(n5650), .Y(n4613) );
  MUX2X1 U5205 ( .B(n4612), .A(n4609), .S(n5727), .Y(n4623) );
  MUX2X1 U5206 ( .B(fifo_array[261]), .A(fifo_array[303]), .S(n5651), .Y(n4617) );
  MUX2X1 U5207 ( .B(fifo_array[177]), .A(fifo_array[219]), .S(n5651), .Y(n4616) );
  MUX2X1 U5208 ( .B(fifo_array[93]), .A(fifo_array[135]), .S(n5651), .Y(n4620)
         );
  MUX2X1 U5209 ( .B(fifo_array[9]), .A(fifo_array[51]), .S(n5651), .Y(n4619)
         );
  MUX2X1 U5210 ( .B(n4618), .A(n4615), .S(n5727), .Y(n4622) );
  MUX2X1 U5211 ( .B(n4621), .A(n4606), .S(n23), .Y(n5593) );
  MUX2X1 U5212 ( .B(fifo_array[1270]), .A(fifo_array[1312]), .S(n5651), .Y(
        n4626) );
  MUX2X1 U5213 ( .B(fifo_array[1186]), .A(fifo_array[1228]), .S(n5651), .Y(
        n4625) );
  MUX2X1 U5214 ( .B(fifo_array[1102]), .A(fifo_array[1144]), .S(n5651), .Y(
        n4629) );
  MUX2X1 U5215 ( .B(fifo_array[1018]), .A(fifo_array[1060]), .S(n5651), .Y(
        n4628) );
  MUX2X1 U5216 ( .B(n4627), .A(n4624), .S(n5727), .Y(n4638) );
  MUX2X1 U5217 ( .B(fifo_array[934]), .A(fifo_array[976]), .S(n5651), .Y(n4632) );
  MUX2X1 U5218 ( .B(fifo_array[850]), .A(fifo_array[892]), .S(n5651), .Y(n4631) );
  MUX2X1 U5219 ( .B(fifo_array[766]), .A(fifo_array[808]), .S(n5651), .Y(n4635) );
  MUX2X1 U5220 ( .B(fifo_array[682]), .A(fifo_array[724]), .S(n5651), .Y(n4634) );
  MUX2X1 U5221 ( .B(n4633), .A(n4630), .S(n5727), .Y(n4637) );
  MUX2X1 U5222 ( .B(fifo_array[598]), .A(fifo_array[640]), .S(n5652), .Y(n4641) );
  MUX2X1 U5223 ( .B(fifo_array[514]), .A(fifo_array[556]), .S(n5652), .Y(n4640) );
  MUX2X1 U5224 ( .B(fifo_array[430]), .A(fifo_array[472]), .S(n5652), .Y(n4644) );
  MUX2X1 U5225 ( .B(fifo_array[346]), .A(fifo_array[388]), .S(n5652), .Y(n4643) );
  MUX2X1 U5226 ( .B(n4642), .A(n4639), .S(n5727), .Y(n4653) );
  MUX2X1 U5227 ( .B(fifo_array[262]), .A(fifo_array[304]), .S(n5652), .Y(n4647) );
  MUX2X1 U5228 ( .B(fifo_array[178]), .A(fifo_array[220]), .S(n5652), .Y(n4646) );
  MUX2X1 U5229 ( .B(fifo_array[94]), .A(fifo_array[136]), .S(n5652), .Y(n4650)
         );
  MUX2X1 U5230 ( .B(fifo_array[10]), .A(fifo_array[52]), .S(n5652), .Y(n4649)
         );
  MUX2X1 U5231 ( .B(n4648), .A(n4645), .S(n5727), .Y(n4652) );
  MUX2X1 U5232 ( .B(n4651), .A(n4636), .S(n23), .Y(n5594) );
  MUX2X1 U5233 ( .B(fifo_array[1271]), .A(fifo_array[1313]), .S(n5652), .Y(
        n4656) );
  MUX2X1 U5234 ( .B(fifo_array[1187]), .A(fifo_array[1229]), .S(n5652), .Y(
        n4655) );
  MUX2X1 U5235 ( .B(fifo_array[1103]), .A(fifo_array[1145]), .S(n5652), .Y(
        n4659) );
  MUX2X1 U5236 ( .B(fifo_array[1019]), .A(fifo_array[1061]), .S(n5652), .Y(
        n4658) );
  MUX2X1 U5237 ( .B(n4657), .A(n4654), .S(n5727), .Y(n4668) );
  MUX2X1 U5238 ( .B(fifo_array[935]), .A(fifo_array[977]), .S(n5653), .Y(n4662) );
  MUX2X1 U5239 ( .B(fifo_array[851]), .A(fifo_array[893]), .S(n5653), .Y(n4661) );
  MUX2X1 U5240 ( .B(fifo_array[767]), .A(fifo_array[809]), .S(n5653), .Y(n4665) );
  MUX2X1 U5241 ( .B(fifo_array[683]), .A(fifo_array[725]), .S(n5653), .Y(n4664) );
  MUX2X1 U5242 ( .B(n4663), .A(n4660), .S(n5727), .Y(n4667) );
  MUX2X1 U5243 ( .B(fifo_array[599]), .A(fifo_array[641]), .S(n5653), .Y(n4671) );
  MUX2X1 U5244 ( .B(fifo_array[515]), .A(fifo_array[557]), .S(n5653), .Y(n4670) );
  MUX2X1 U5245 ( .B(fifo_array[431]), .A(fifo_array[473]), .S(n5653), .Y(n4674) );
  MUX2X1 U5246 ( .B(fifo_array[347]), .A(fifo_array[389]), .S(n5653), .Y(n4673) );
  MUX2X1 U5247 ( .B(n4672), .A(n4669), .S(n5727), .Y(n4683) );
  MUX2X1 U5248 ( .B(fifo_array[263]), .A(fifo_array[305]), .S(n5653), .Y(n4677) );
  MUX2X1 U5249 ( .B(fifo_array[179]), .A(fifo_array[221]), .S(n5653), .Y(n4676) );
  MUX2X1 U5250 ( .B(fifo_array[95]), .A(fifo_array[137]), .S(n5653), .Y(n4680)
         );
  MUX2X1 U5251 ( .B(fifo_array[11]), .A(fifo_array[53]), .S(n5653), .Y(n4679)
         );
  MUX2X1 U5252 ( .B(n4678), .A(n4675), .S(n5727), .Y(n4682) );
  MUX2X1 U5253 ( .B(n4681), .A(n4666), .S(n23), .Y(n5595) );
  MUX2X1 U5254 ( .B(fifo_array[1272]), .A(fifo_array[1314]), .S(n5654), .Y(
        n4686) );
  MUX2X1 U5255 ( .B(fifo_array[1188]), .A(fifo_array[1230]), .S(n5654), .Y(
        n4685) );
  MUX2X1 U5256 ( .B(fifo_array[1104]), .A(fifo_array[1146]), .S(n5654), .Y(
        n4689) );
  MUX2X1 U5257 ( .B(fifo_array[1020]), .A(fifo_array[1062]), .S(n5654), .Y(
        n4688) );
  MUX2X1 U5258 ( .B(n4687), .A(n4684), .S(n5728), .Y(n4698) );
  MUX2X1 U5259 ( .B(fifo_array[936]), .A(fifo_array[978]), .S(n5654), .Y(n4692) );
  MUX2X1 U5260 ( .B(fifo_array[852]), .A(fifo_array[894]), .S(n5654), .Y(n4691) );
  MUX2X1 U5261 ( .B(fifo_array[768]), .A(fifo_array[810]), .S(n5654), .Y(n4695) );
  MUX2X1 U5262 ( .B(fifo_array[684]), .A(fifo_array[726]), .S(n5654), .Y(n4694) );
  MUX2X1 U5263 ( .B(n4693), .A(n4690), .S(n5728), .Y(n4697) );
  MUX2X1 U5264 ( .B(fifo_array[600]), .A(fifo_array[642]), .S(n5654), .Y(n4701) );
  MUX2X1 U5265 ( .B(fifo_array[516]), .A(fifo_array[558]), .S(n5654), .Y(n4700) );
  MUX2X1 U5266 ( .B(fifo_array[432]), .A(fifo_array[474]), .S(n5654), .Y(n4704) );
  MUX2X1 U5267 ( .B(fifo_array[348]), .A(fifo_array[390]), .S(n5654), .Y(n4703) );
  MUX2X1 U5268 ( .B(n4702), .A(n4699), .S(n5728), .Y(n4713) );
  MUX2X1 U5269 ( .B(fifo_array[264]), .A(fifo_array[306]), .S(n5655), .Y(n4707) );
  MUX2X1 U5270 ( .B(fifo_array[180]), .A(fifo_array[222]), .S(n5655), .Y(n4706) );
  MUX2X1 U5271 ( .B(fifo_array[96]), .A(fifo_array[138]), .S(n5655), .Y(n4710)
         );
  MUX2X1 U5272 ( .B(fifo_array[12]), .A(fifo_array[54]), .S(n5655), .Y(n4709)
         );
  MUX2X1 U5273 ( .B(n4708), .A(n4705), .S(n5728), .Y(n4712) );
  MUX2X1 U5274 ( .B(n4711), .A(n4696), .S(n23), .Y(n5596) );
  MUX2X1 U5275 ( .B(fifo_array[1273]), .A(fifo_array[1315]), .S(n5655), .Y(
        n4716) );
  MUX2X1 U5276 ( .B(fifo_array[1189]), .A(fifo_array[1231]), .S(n5655), .Y(
        n4715) );
  MUX2X1 U5277 ( .B(fifo_array[1105]), .A(fifo_array[1147]), .S(n5655), .Y(
        n4719) );
  MUX2X1 U5278 ( .B(fifo_array[1021]), .A(fifo_array[1063]), .S(n5655), .Y(
        n4718) );
  MUX2X1 U5279 ( .B(n4717), .A(n4714), .S(n5728), .Y(n4728) );
  MUX2X1 U5280 ( .B(fifo_array[937]), .A(fifo_array[979]), .S(n5655), .Y(n4722) );
  MUX2X1 U5281 ( .B(fifo_array[853]), .A(fifo_array[895]), .S(n5655), .Y(n4721) );
  MUX2X1 U5282 ( .B(fifo_array[769]), .A(fifo_array[811]), .S(n5655), .Y(n4725) );
  MUX2X1 U5283 ( .B(fifo_array[685]), .A(fifo_array[727]), .S(n5655), .Y(n4724) );
  MUX2X1 U5284 ( .B(n4723), .A(n4720), .S(n5728), .Y(n4727) );
  MUX2X1 U5285 ( .B(fifo_array[601]), .A(fifo_array[643]), .S(n5656), .Y(n4731) );
  MUX2X1 U5286 ( .B(fifo_array[517]), .A(fifo_array[559]), .S(n5656), .Y(n4730) );
  MUX2X1 U5287 ( .B(fifo_array[433]), .A(fifo_array[475]), .S(n5656), .Y(n4734) );
  MUX2X1 U5288 ( .B(fifo_array[349]), .A(fifo_array[391]), .S(n5656), .Y(n4733) );
  MUX2X1 U5289 ( .B(n4732), .A(n4729), .S(n5728), .Y(n4743) );
  MUX2X1 U5290 ( .B(fifo_array[265]), .A(fifo_array[307]), .S(n5656), .Y(n4737) );
  MUX2X1 U5291 ( .B(fifo_array[181]), .A(fifo_array[223]), .S(n5656), .Y(n4736) );
  MUX2X1 U5292 ( .B(fifo_array[97]), .A(fifo_array[139]), .S(n5656), .Y(n4740)
         );
  MUX2X1 U5293 ( .B(fifo_array[13]), .A(fifo_array[55]), .S(n5656), .Y(n4739)
         );
  MUX2X1 U5294 ( .B(n4738), .A(n4735), .S(n5728), .Y(n4742) );
  MUX2X1 U5295 ( .B(n4741), .A(n4726), .S(n23), .Y(n5597) );
  MUX2X1 U5296 ( .B(fifo_array[1274]), .A(fifo_array[1316]), .S(n5656), .Y(
        n4746) );
  MUX2X1 U5297 ( .B(fifo_array[1190]), .A(fifo_array[1232]), .S(n5656), .Y(
        n4745) );
  MUX2X1 U5298 ( .B(fifo_array[1106]), .A(fifo_array[1148]), .S(n5656), .Y(
        n4749) );
  MUX2X1 U5299 ( .B(fifo_array[1022]), .A(fifo_array[1064]), .S(n5656), .Y(
        n4748) );
  MUX2X1 U5300 ( .B(n4747), .A(n4744), .S(n5728), .Y(n4758) );
  MUX2X1 U5301 ( .B(fifo_array[938]), .A(fifo_array[980]), .S(n5657), .Y(n4752) );
  MUX2X1 U5302 ( .B(fifo_array[854]), .A(fifo_array[896]), .S(n5657), .Y(n4751) );
  MUX2X1 U5303 ( .B(fifo_array[770]), .A(fifo_array[812]), .S(n5657), .Y(n4755) );
  MUX2X1 U5304 ( .B(fifo_array[686]), .A(fifo_array[728]), .S(n5657), .Y(n4754) );
  MUX2X1 U5305 ( .B(n4753), .A(n4750), .S(n5728), .Y(n4757) );
  MUX2X1 U5306 ( .B(fifo_array[602]), .A(fifo_array[644]), .S(n5657), .Y(n4761) );
  MUX2X1 U5307 ( .B(fifo_array[518]), .A(fifo_array[560]), .S(n5657), .Y(n4760) );
  MUX2X1 U5308 ( .B(fifo_array[434]), .A(fifo_array[476]), .S(n5657), .Y(n4764) );
  MUX2X1 U5309 ( .B(fifo_array[350]), .A(fifo_array[392]), .S(n5657), .Y(n4763) );
  MUX2X1 U5310 ( .B(n4762), .A(n4759), .S(n5728), .Y(n4773) );
  MUX2X1 U5311 ( .B(fifo_array[266]), .A(fifo_array[308]), .S(n5657), .Y(n4767) );
  MUX2X1 U5312 ( .B(fifo_array[182]), .A(fifo_array[224]), .S(n5657), .Y(n4766) );
  MUX2X1 U5313 ( .B(fifo_array[98]), .A(fifo_array[140]), .S(n5657), .Y(n4770)
         );
  MUX2X1 U5314 ( .B(fifo_array[14]), .A(fifo_array[56]), .S(n5657), .Y(n4769)
         );
  MUX2X1 U5315 ( .B(n4768), .A(n4765), .S(n5728), .Y(n4772) );
  MUX2X1 U5316 ( .B(n4771), .A(n4756), .S(n23), .Y(n5598) );
  MUX2X1 U5317 ( .B(fifo_array[1275]), .A(fifo_array[1317]), .S(n5658), .Y(
        n4776) );
  MUX2X1 U5318 ( .B(fifo_array[1191]), .A(fifo_array[1233]), .S(n5658), .Y(
        n4775) );
  MUX2X1 U5319 ( .B(fifo_array[1107]), .A(fifo_array[1149]), .S(n5658), .Y(
        n4779) );
  MUX2X1 U5320 ( .B(fifo_array[1023]), .A(fifo_array[1065]), .S(n5658), .Y(
        n4778) );
  MUX2X1 U5321 ( .B(n4777), .A(n4774), .S(n5729), .Y(n4788) );
  MUX2X1 U5322 ( .B(fifo_array[939]), .A(fifo_array[981]), .S(n5658), .Y(n4782) );
  MUX2X1 U5323 ( .B(fifo_array[855]), .A(fifo_array[897]), .S(n5658), .Y(n4781) );
  MUX2X1 U5324 ( .B(fifo_array[771]), .A(fifo_array[813]), .S(n5658), .Y(n4785) );
  MUX2X1 U5325 ( .B(fifo_array[687]), .A(fifo_array[729]), .S(n5658), .Y(n4784) );
  MUX2X1 U5326 ( .B(n4783), .A(n4780), .S(n5729), .Y(n4787) );
  MUX2X1 U5327 ( .B(fifo_array[603]), .A(fifo_array[645]), .S(n5658), .Y(n4791) );
  MUX2X1 U5328 ( .B(fifo_array[519]), .A(fifo_array[561]), .S(n5658), .Y(n4790) );
  MUX2X1 U5329 ( .B(fifo_array[435]), .A(fifo_array[477]), .S(n5658), .Y(n4794) );
  MUX2X1 U5330 ( .B(fifo_array[351]), .A(fifo_array[393]), .S(n5658), .Y(n4793) );
  MUX2X1 U5331 ( .B(n4792), .A(n4789), .S(n5729), .Y(n4803) );
  MUX2X1 U5332 ( .B(fifo_array[267]), .A(fifo_array[309]), .S(n5659), .Y(n4797) );
  MUX2X1 U5333 ( .B(fifo_array[183]), .A(fifo_array[225]), .S(n5659), .Y(n4796) );
  MUX2X1 U5334 ( .B(fifo_array[99]), .A(fifo_array[141]), .S(n5659), .Y(n4800)
         );
  MUX2X1 U5335 ( .B(fifo_array[15]), .A(fifo_array[57]), .S(n5659), .Y(n4799)
         );
  MUX2X1 U5336 ( .B(n4798), .A(n4795), .S(n5729), .Y(n4802) );
  MUX2X1 U5337 ( .B(n4801), .A(n4786), .S(n23), .Y(n5599) );
  MUX2X1 U5338 ( .B(fifo_array[1276]), .A(fifo_array[1318]), .S(n5659), .Y(
        n4806) );
  MUX2X1 U5339 ( .B(fifo_array[1192]), .A(fifo_array[1234]), .S(n5659), .Y(
        n4805) );
  MUX2X1 U5340 ( .B(fifo_array[1108]), .A(fifo_array[1150]), .S(n5659), .Y(
        n4809) );
  MUX2X1 U5341 ( .B(fifo_array[1024]), .A(fifo_array[1066]), .S(n5659), .Y(
        n4808) );
  MUX2X1 U5342 ( .B(n4807), .A(n4804), .S(n5729), .Y(n4818) );
  MUX2X1 U5343 ( .B(fifo_array[940]), .A(fifo_array[982]), .S(n5659), .Y(n4812) );
  MUX2X1 U5344 ( .B(fifo_array[856]), .A(fifo_array[898]), .S(n5659), .Y(n4811) );
  MUX2X1 U5345 ( .B(fifo_array[772]), .A(fifo_array[814]), .S(n5659), .Y(n4815) );
  MUX2X1 U5346 ( .B(fifo_array[688]), .A(fifo_array[730]), .S(n5659), .Y(n4814) );
  MUX2X1 U5347 ( .B(n4813), .A(n4810), .S(n5729), .Y(n4817) );
  MUX2X1 U5348 ( .B(fifo_array[604]), .A(fifo_array[646]), .S(n5660), .Y(n4821) );
  MUX2X1 U5349 ( .B(fifo_array[520]), .A(fifo_array[562]), .S(n5660), .Y(n4820) );
  MUX2X1 U5350 ( .B(fifo_array[436]), .A(fifo_array[478]), .S(n5660), .Y(n4824) );
  MUX2X1 U5351 ( .B(fifo_array[352]), .A(fifo_array[394]), .S(n5660), .Y(n4823) );
  MUX2X1 U5352 ( .B(n4822), .A(n4819), .S(n5729), .Y(n4833) );
  MUX2X1 U5353 ( .B(fifo_array[268]), .A(fifo_array[310]), .S(n5660), .Y(n4827) );
  MUX2X1 U5354 ( .B(fifo_array[184]), .A(fifo_array[226]), .S(n5660), .Y(n4826) );
  MUX2X1 U5355 ( .B(fifo_array[100]), .A(fifo_array[142]), .S(n5660), .Y(n4830) );
  MUX2X1 U5356 ( .B(fifo_array[16]), .A(fifo_array[58]), .S(n5660), .Y(n4829)
         );
  MUX2X1 U5357 ( .B(n4828), .A(n4825), .S(n5729), .Y(n4832) );
  MUX2X1 U5358 ( .B(n4831), .A(n4816), .S(n23), .Y(n5600) );
  MUX2X1 U5359 ( .B(fifo_array[1277]), .A(fifo_array[1319]), .S(n5660), .Y(
        n4836) );
  MUX2X1 U5360 ( .B(fifo_array[1193]), .A(fifo_array[1235]), .S(n5660), .Y(
        n4835) );
  MUX2X1 U5361 ( .B(fifo_array[1109]), .A(fifo_array[1151]), .S(n5660), .Y(
        n4839) );
  MUX2X1 U5362 ( .B(fifo_array[1025]), .A(fifo_array[1067]), .S(n5660), .Y(
        n4838) );
  MUX2X1 U5363 ( .B(n4837), .A(n4834), .S(n5729), .Y(n4848) );
  MUX2X1 U5364 ( .B(fifo_array[941]), .A(fifo_array[983]), .S(n5661), .Y(n4842) );
  MUX2X1 U5365 ( .B(fifo_array[857]), .A(fifo_array[899]), .S(n5661), .Y(n4841) );
  MUX2X1 U5366 ( .B(fifo_array[773]), .A(fifo_array[815]), .S(n5661), .Y(n4845) );
  MUX2X1 U5367 ( .B(fifo_array[689]), .A(fifo_array[731]), .S(n5661), .Y(n4844) );
  MUX2X1 U5368 ( .B(n4843), .A(n4840), .S(n5729), .Y(n4847) );
  MUX2X1 U5369 ( .B(fifo_array[605]), .A(fifo_array[647]), .S(n5661), .Y(n4851) );
  MUX2X1 U5370 ( .B(fifo_array[521]), .A(fifo_array[563]), .S(n5661), .Y(n4850) );
  MUX2X1 U5371 ( .B(fifo_array[437]), .A(fifo_array[479]), .S(n5661), .Y(n4854) );
  MUX2X1 U5372 ( .B(fifo_array[353]), .A(fifo_array[395]), .S(n5661), .Y(n4853) );
  MUX2X1 U5373 ( .B(n4852), .A(n4849), .S(n5729), .Y(n4863) );
  MUX2X1 U5374 ( .B(fifo_array[269]), .A(fifo_array[311]), .S(n5661), .Y(n4857) );
  MUX2X1 U5375 ( .B(fifo_array[185]), .A(fifo_array[227]), .S(n5661), .Y(n4856) );
  MUX2X1 U5376 ( .B(fifo_array[101]), .A(fifo_array[143]), .S(n5661), .Y(n4860) );
  MUX2X1 U5377 ( .B(fifo_array[17]), .A(fifo_array[59]), .S(n5661), .Y(n4859)
         );
  MUX2X1 U5378 ( .B(n4858), .A(n4855), .S(n5729), .Y(n4862) );
  MUX2X1 U5379 ( .B(n4861), .A(n4846), .S(n23), .Y(n5601) );
  MUX2X1 U5380 ( .B(fifo_array[1278]), .A(fifo_array[1320]), .S(n5662), .Y(
        n4866) );
  MUX2X1 U5381 ( .B(fifo_array[1194]), .A(fifo_array[1236]), .S(n5662), .Y(
        n4865) );
  MUX2X1 U5382 ( .B(fifo_array[1110]), .A(fifo_array[1152]), .S(n5662), .Y(
        n4869) );
  MUX2X1 U5383 ( .B(fifo_array[1026]), .A(fifo_array[1068]), .S(n5662), .Y(
        n4868) );
  MUX2X1 U5384 ( .B(n4867), .A(n4864), .S(n5725), .Y(n4878) );
  MUX2X1 U5385 ( .B(fifo_array[942]), .A(fifo_array[984]), .S(n5662), .Y(n4872) );
  MUX2X1 U5386 ( .B(fifo_array[858]), .A(fifo_array[900]), .S(n5662), .Y(n4871) );
  MUX2X1 U5387 ( .B(fifo_array[774]), .A(fifo_array[816]), .S(n5662), .Y(n4875) );
  MUX2X1 U5388 ( .B(fifo_array[690]), .A(fifo_array[732]), .S(n5662), .Y(n4874) );
  MUX2X1 U5389 ( .B(n4873), .A(n4870), .S(n21), .Y(n4877) );
  MUX2X1 U5390 ( .B(fifo_array[606]), .A(fifo_array[648]), .S(n5662), .Y(n4881) );
  MUX2X1 U5391 ( .B(fifo_array[522]), .A(fifo_array[564]), .S(n5662), .Y(n4880) );
  MUX2X1 U5392 ( .B(fifo_array[438]), .A(fifo_array[480]), .S(n5662), .Y(n4884) );
  MUX2X1 U5393 ( .B(fifo_array[354]), .A(fifo_array[396]), .S(n5662), .Y(n4883) );
  MUX2X1 U5394 ( .B(n4882), .A(n4879), .S(n5725), .Y(n4893) );
  MUX2X1 U5395 ( .B(fifo_array[270]), .A(fifo_array[312]), .S(n5663), .Y(n4887) );
  MUX2X1 U5396 ( .B(fifo_array[186]), .A(fifo_array[228]), .S(n5663), .Y(n4886) );
  MUX2X1 U5397 ( .B(fifo_array[102]), .A(fifo_array[144]), .S(n5663), .Y(n4890) );
  MUX2X1 U5398 ( .B(fifo_array[18]), .A(fifo_array[60]), .S(n5663), .Y(n4889)
         );
  MUX2X1 U5399 ( .B(n4888), .A(n4885), .S(n5724), .Y(n4892) );
  MUX2X1 U5400 ( .B(n4891), .A(n4876), .S(n23), .Y(n5602) );
  MUX2X1 U5401 ( .B(fifo_array[1279]), .A(fifo_array[1321]), .S(n5663), .Y(
        n4896) );
  MUX2X1 U5402 ( .B(fifo_array[1195]), .A(fifo_array[1237]), .S(n5663), .Y(
        n4895) );
  MUX2X1 U5403 ( .B(fifo_array[1111]), .A(fifo_array[1153]), .S(n5663), .Y(
        n4899) );
  MUX2X1 U5404 ( .B(fifo_array[1027]), .A(fifo_array[1069]), .S(n5663), .Y(
        n4898) );
  MUX2X1 U5405 ( .B(n4897), .A(n4894), .S(n5724), .Y(n4908) );
  MUX2X1 U5406 ( .B(fifo_array[943]), .A(fifo_array[985]), .S(n5663), .Y(n4902) );
  MUX2X1 U5407 ( .B(fifo_array[859]), .A(fifo_array[901]), .S(n5663), .Y(n4901) );
  MUX2X1 U5408 ( .B(fifo_array[775]), .A(fifo_array[817]), .S(n5663), .Y(n4905) );
  MUX2X1 U5409 ( .B(fifo_array[691]), .A(fifo_array[733]), .S(n5663), .Y(n4904) );
  MUX2X1 U5410 ( .B(n4903), .A(n4900), .S(n21), .Y(n4907) );
  MUX2X1 U5411 ( .B(fifo_array[607]), .A(fifo_array[649]), .S(n5664), .Y(n4911) );
  MUX2X1 U5412 ( .B(fifo_array[523]), .A(fifo_array[565]), .S(n5664), .Y(n4910) );
  MUX2X1 U5413 ( .B(fifo_array[439]), .A(fifo_array[481]), .S(n5664), .Y(n4914) );
  MUX2X1 U5414 ( .B(fifo_array[355]), .A(fifo_array[397]), .S(n5664), .Y(n4913) );
  MUX2X1 U5415 ( .B(n4912), .A(n4909), .S(n5724), .Y(n4923) );
  MUX2X1 U5416 ( .B(fifo_array[271]), .A(fifo_array[313]), .S(n5664), .Y(n4917) );
  MUX2X1 U5417 ( .B(fifo_array[187]), .A(fifo_array[229]), .S(n5664), .Y(n4916) );
  MUX2X1 U5418 ( .B(fifo_array[103]), .A(fifo_array[145]), .S(n5664), .Y(n4920) );
  MUX2X1 U5419 ( .B(fifo_array[19]), .A(fifo_array[61]), .S(n5664), .Y(n4919)
         );
  MUX2X1 U5420 ( .B(n4918), .A(n4915), .S(n5725), .Y(n4922) );
  MUX2X1 U5421 ( .B(n4921), .A(n4906), .S(n23), .Y(n5603) );
  MUX2X1 U5422 ( .B(fifo_array[1280]), .A(fifo_array[1322]), .S(n5664), .Y(
        n4926) );
  MUX2X1 U5423 ( .B(fifo_array[1196]), .A(fifo_array[1238]), .S(n5664), .Y(
        n4925) );
  MUX2X1 U5424 ( .B(fifo_array[1112]), .A(fifo_array[1154]), .S(n5664), .Y(
        n4929) );
  MUX2X1 U5425 ( .B(fifo_array[1028]), .A(fifo_array[1070]), .S(n5664), .Y(
        n4928) );
  MUX2X1 U5426 ( .B(n4927), .A(n4924), .S(n21), .Y(n4938) );
  MUX2X1 U5427 ( .B(fifo_array[944]), .A(fifo_array[986]), .S(n5665), .Y(n4932) );
  MUX2X1 U5428 ( .B(fifo_array[860]), .A(fifo_array[902]), .S(n5665), .Y(n4931) );
  MUX2X1 U5429 ( .B(fifo_array[776]), .A(fifo_array[818]), .S(n5665), .Y(n4935) );
  MUX2X1 U5430 ( .B(fifo_array[692]), .A(fifo_array[734]), .S(n5665), .Y(n4934) );
  MUX2X1 U5431 ( .B(n4933), .A(n4930), .S(n21), .Y(n4937) );
  MUX2X1 U5432 ( .B(fifo_array[608]), .A(fifo_array[650]), .S(n5665), .Y(n4941) );
  MUX2X1 U5433 ( .B(fifo_array[524]), .A(fifo_array[566]), .S(n5665), .Y(n4940) );
  MUX2X1 U5434 ( .B(fifo_array[440]), .A(fifo_array[482]), .S(n5665), .Y(n4944) );
  MUX2X1 U5435 ( .B(fifo_array[356]), .A(fifo_array[398]), .S(n5665), .Y(n4943) );
  MUX2X1 U5436 ( .B(n4942), .A(n4939), .S(n5725), .Y(n4953) );
  MUX2X1 U5437 ( .B(fifo_array[272]), .A(fifo_array[314]), .S(n5665), .Y(n4947) );
  MUX2X1 U5438 ( .B(fifo_array[188]), .A(fifo_array[230]), .S(n5665), .Y(n4946) );
  MUX2X1 U5439 ( .B(fifo_array[104]), .A(fifo_array[146]), .S(n5665), .Y(n4950) );
  MUX2X1 U5440 ( .B(fifo_array[20]), .A(fifo_array[62]), .S(n5665), .Y(n4949)
         );
  MUX2X1 U5441 ( .B(n4948), .A(n4945), .S(n5724), .Y(n4952) );
  MUX2X1 U5442 ( .B(n4951), .A(n4936), .S(n23), .Y(n5604) );
  MUX2X1 U5443 ( .B(fifo_array[1281]), .A(fifo_array[1323]), .S(n5666), .Y(
        n4956) );
  MUX2X1 U5444 ( .B(fifo_array[1197]), .A(fifo_array[1239]), .S(n5666), .Y(
        n4955) );
  MUX2X1 U5445 ( .B(fifo_array[1113]), .A(fifo_array[1155]), .S(n5666), .Y(
        n4959) );
  MUX2X1 U5446 ( .B(fifo_array[1029]), .A(fifo_array[1071]), .S(n5666), .Y(
        n4958) );
  MUX2X1 U5447 ( .B(n4957), .A(n4954), .S(n21), .Y(n4968) );
  MUX2X1 U5448 ( .B(fifo_array[945]), .A(fifo_array[987]), .S(n5666), .Y(n4962) );
  MUX2X1 U5449 ( .B(fifo_array[861]), .A(fifo_array[903]), .S(n5666), .Y(n4961) );
  MUX2X1 U5450 ( .B(fifo_array[777]), .A(fifo_array[819]), .S(n5666), .Y(n4965) );
  MUX2X1 U5451 ( .B(fifo_array[693]), .A(fifo_array[735]), .S(n5666), .Y(n4964) );
  MUX2X1 U5452 ( .B(n4963), .A(n4960), .S(n21), .Y(n4967) );
  MUX2X1 U5453 ( .B(fifo_array[609]), .A(fifo_array[651]), .S(n5666), .Y(n4971) );
  MUX2X1 U5454 ( .B(fifo_array[525]), .A(fifo_array[567]), .S(n5666), .Y(n4970) );
  MUX2X1 U5455 ( .B(fifo_array[441]), .A(fifo_array[483]), .S(n5666), .Y(n4974) );
  MUX2X1 U5456 ( .B(fifo_array[357]), .A(fifo_array[399]), .S(n5666), .Y(n4973) );
  MUX2X1 U5457 ( .B(n4972), .A(n4969), .S(n5728), .Y(n4983) );
  MUX2X1 U5458 ( .B(fifo_array[273]), .A(fifo_array[315]), .S(n5667), .Y(n4977) );
  MUX2X1 U5459 ( .B(fifo_array[189]), .A(fifo_array[231]), .S(n5667), .Y(n4976) );
  MUX2X1 U5460 ( .B(fifo_array[105]), .A(fifo_array[147]), .S(n5667), .Y(n4980) );
  MUX2X1 U5461 ( .B(fifo_array[21]), .A(fifo_array[63]), .S(n5667), .Y(n4979)
         );
  MUX2X1 U5462 ( .B(n4978), .A(n4975), .S(n5727), .Y(n4982) );
  MUX2X1 U5463 ( .B(n4981), .A(n4966), .S(n23), .Y(n5605) );
  MUX2X1 U5464 ( .B(fifo_array[1282]), .A(fifo_array[1324]), .S(n5667), .Y(
        n4986) );
  MUX2X1 U5465 ( .B(fifo_array[1198]), .A(fifo_array[1240]), .S(n5667), .Y(
        n4985) );
  MUX2X1 U5466 ( .B(fifo_array[1114]), .A(fifo_array[1156]), .S(n5667), .Y(
        n4989) );
  MUX2X1 U5467 ( .B(fifo_array[1030]), .A(fifo_array[1072]), .S(n5667), .Y(
        n4988) );
  MUX2X1 U5468 ( .B(n4987), .A(n4984), .S(n21), .Y(n4998) );
  MUX2X1 U5469 ( .B(fifo_array[946]), .A(fifo_array[988]), .S(n5667), .Y(n4992) );
  MUX2X1 U5470 ( .B(fifo_array[862]), .A(fifo_array[904]), .S(n5667), .Y(n4991) );
  MUX2X1 U5471 ( .B(fifo_array[778]), .A(fifo_array[820]), .S(n5667), .Y(n4995) );
  MUX2X1 U5472 ( .B(fifo_array[694]), .A(fifo_array[736]), .S(n5667), .Y(n4994) );
  MUX2X1 U5473 ( .B(n4993), .A(n4990), .S(n21), .Y(n4997) );
  MUX2X1 U5474 ( .B(fifo_array[610]), .A(fifo_array[652]), .S(n5668), .Y(n5001) );
  MUX2X1 U5475 ( .B(fifo_array[526]), .A(fifo_array[568]), .S(n5668), .Y(n5000) );
  MUX2X1 U5476 ( .B(fifo_array[442]), .A(fifo_array[484]), .S(n5668), .Y(n5004) );
  MUX2X1 U5477 ( .B(fifo_array[358]), .A(fifo_array[400]), .S(n5668), .Y(n5003) );
  MUX2X1 U5478 ( .B(n5002), .A(n4999), .S(n5728), .Y(n5013) );
  MUX2X1 U5479 ( .B(fifo_array[274]), .A(fifo_array[316]), .S(n5668), .Y(n5007) );
  MUX2X1 U5480 ( .B(fifo_array[190]), .A(fifo_array[232]), .S(n5668), .Y(n5006) );
  MUX2X1 U5481 ( .B(fifo_array[106]), .A(fifo_array[148]), .S(n5668), .Y(n5010) );
  MUX2X1 U5482 ( .B(fifo_array[22]), .A(fifo_array[64]), .S(n5668), .Y(n5009)
         );
  MUX2X1 U5483 ( .B(n5008), .A(n5005), .S(n21), .Y(n5012) );
  MUX2X1 U5484 ( .B(n5011), .A(n4996), .S(n23), .Y(n5606) );
  MUX2X1 U5485 ( .B(fifo_array[1283]), .A(fifo_array[1325]), .S(n5668), .Y(
        n5016) );
  MUX2X1 U5486 ( .B(fifo_array[1199]), .A(fifo_array[1241]), .S(n5668), .Y(
        n5015) );
  MUX2X1 U5487 ( .B(fifo_array[1115]), .A(fifo_array[1157]), .S(n5668), .Y(
        n5019) );
  MUX2X1 U5488 ( .B(fifo_array[1031]), .A(fifo_array[1073]), .S(n5668), .Y(
        n5018) );
  MUX2X1 U5489 ( .B(n5017), .A(n5014), .S(n21), .Y(n5028) );
  MUX2X1 U5490 ( .B(fifo_array[947]), .A(fifo_array[989]), .S(n5669), .Y(n5022) );
  MUX2X1 U5491 ( .B(fifo_array[863]), .A(fifo_array[905]), .S(n5669), .Y(n5021) );
  MUX2X1 U5492 ( .B(fifo_array[779]), .A(fifo_array[821]), .S(n5669), .Y(n5025) );
  MUX2X1 U5493 ( .B(fifo_array[695]), .A(fifo_array[737]), .S(n5669), .Y(n5024) );
  MUX2X1 U5494 ( .B(n5023), .A(n5020), .S(n21), .Y(n5027) );
  MUX2X1 U5495 ( .B(fifo_array[611]), .A(fifo_array[653]), .S(n5669), .Y(n5031) );
  MUX2X1 U5496 ( .B(fifo_array[527]), .A(fifo_array[569]), .S(n5669), .Y(n5030) );
  MUX2X1 U5497 ( .B(fifo_array[443]), .A(fifo_array[485]), .S(n5669), .Y(n5034) );
  MUX2X1 U5498 ( .B(fifo_array[359]), .A(fifo_array[401]), .S(n5669), .Y(n5033) );
  MUX2X1 U5499 ( .B(n5032), .A(n5029), .S(n5729), .Y(n5043) );
  MUX2X1 U5500 ( .B(fifo_array[275]), .A(fifo_array[317]), .S(n5669), .Y(n5037) );
  MUX2X1 U5501 ( .B(fifo_array[191]), .A(fifo_array[233]), .S(n5669), .Y(n5036) );
  MUX2X1 U5502 ( .B(fifo_array[107]), .A(fifo_array[149]), .S(n5669), .Y(n5040) );
  MUX2X1 U5503 ( .B(fifo_array[23]), .A(fifo_array[65]), .S(n5669), .Y(n5039)
         );
  MUX2X1 U5504 ( .B(n5038), .A(n5035), .S(n5726), .Y(n5042) );
  MUX2X1 U5505 ( .B(n5041), .A(n5026), .S(n23), .Y(n5607) );
  MUX2X1 U5506 ( .B(fifo_array[1284]), .A(fifo_array[1326]), .S(n5670), .Y(
        n5046) );
  MUX2X1 U5507 ( .B(fifo_array[1200]), .A(fifo_array[1242]), .S(n5670), .Y(
        n5045) );
  MUX2X1 U5508 ( .B(fifo_array[1116]), .A(fifo_array[1158]), .S(n5670), .Y(
        n5049) );
  MUX2X1 U5509 ( .B(fifo_array[1032]), .A(fifo_array[1074]), .S(n5670), .Y(
        n5048) );
  MUX2X1 U5510 ( .B(n5047), .A(n5044), .S(n5727), .Y(n5058) );
  MUX2X1 U5511 ( .B(fifo_array[948]), .A(fifo_array[990]), .S(n5670), .Y(n5052) );
  MUX2X1 U5512 ( .B(fifo_array[864]), .A(fifo_array[906]), .S(n5670), .Y(n5051) );
  MUX2X1 U5513 ( .B(fifo_array[780]), .A(fifo_array[822]), .S(n5670), .Y(n5055) );
  MUX2X1 U5514 ( .B(fifo_array[696]), .A(fifo_array[738]), .S(n5670), .Y(n5054) );
  MUX2X1 U5515 ( .B(n5053), .A(n5050), .S(n5729), .Y(n5057) );
  MUX2X1 U5516 ( .B(fifo_array[612]), .A(fifo_array[654]), .S(n5670), .Y(n5061) );
  MUX2X1 U5517 ( .B(fifo_array[528]), .A(fifo_array[570]), .S(n5670), .Y(n5060) );
  MUX2X1 U5518 ( .B(fifo_array[444]), .A(fifo_array[486]), .S(n5670), .Y(n5064) );
  MUX2X1 U5519 ( .B(fifo_array[360]), .A(fifo_array[402]), .S(n5670), .Y(n5063) );
  MUX2X1 U5520 ( .B(n5062), .A(n5059), .S(n5729), .Y(n5073) );
  MUX2X1 U5521 ( .B(fifo_array[276]), .A(fifo_array[318]), .S(n5671), .Y(n5067) );
  MUX2X1 U5522 ( .B(fifo_array[192]), .A(fifo_array[234]), .S(n5671), .Y(n5066) );
  MUX2X1 U5523 ( .B(fifo_array[108]), .A(fifo_array[150]), .S(n5671), .Y(n5070) );
  MUX2X1 U5524 ( .B(fifo_array[24]), .A(fifo_array[66]), .S(n5671), .Y(n5069)
         );
  MUX2X1 U5525 ( .B(n5068), .A(n5065), .S(n5726), .Y(n5072) );
  MUX2X1 U5526 ( .B(n5071), .A(n5056), .S(n23), .Y(n5608) );
  MUX2X1 U5527 ( .B(fifo_array[1285]), .A(fifo_array[1327]), .S(n5671), .Y(
        n5076) );
  MUX2X1 U5528 ( .B(fifo_array[1201]), .A(fifo_array[1243]), .S(n5671), .Y(
        n5075) );
  MUX2X1 U5529 ( .B(fifo_array[1117]), .A(fifo_array[1159]), .S(n5671), .Y(
        n5079) );
  MUX2X1 U5530 ( .B(fifo_array[1033]), .A(fifo_array[1075]), .S(n5671), .Y(
        n5078) );
  MUX2X1 U5531 ( .B(n5077), .A(n5074), .S(n21), .Y(n5088) );
  MUX2X1 U5532 ( .B(fifo_array[949]), .A(fifo_array[991]), .S(n5671), .Y(n5082) );
  MUX2X1 U5533 ( .B(fifo_array[865]), .A(fifo_array[907]), .S(n5671), .Y(n5081) );
  MUX2X1 U5534 ( .B(fifo_array[781]), .A(fifo_array[823]), .S(n5671), .Y(n5085) );
  MUX2X1 U5535 ( .B(fifo_array[697]), .A(fifo_array[739]), .S(n5671), .Y(n5084) );
  MUX2X1 U5536 ( .B(n5083), .A(n5080), .S(n5726), .Y(n5087) );
  MUX2X1 U5537 ( .B(fifo_array[613]), .A(fifo_array[655]), .S(n5672), .Y(n5091) );
  MUX2X1 U5538 ( .B(fifo_array[529]), .A(fifo_array[571]), .S(n5672), .Y(n5090) );
  MUX2X1 U5539 ( .B(fifo_array[445]), .A(fifo_array[487]), .S(n5672), .Y(n5094) );
  MUX2X1 U5540 ( .B(fifo_array[361]), .A(fifo_array[403]), .S(n5672), .Y(n5093) );
  MUX2X1 U5541 ( .B(n5092), .A(n5089), .S(n5728), .Y(n5103) );
  MUX2X1 U5542 ( .B(fifo_array[277]), .A(fifo_array[319]), .S(n5672), .Y(n5097) );
  MUX2X1 U5543 ( .B(fifo_array[193]), .A(fifo_array[235]), .S(n5672), .Y(n5096) );
  MUX2X1 U5544 ( .B(fifo_array[109]), .A(fifo_array[151]), .S(n5672), .Y(n5100) );
  MUX2X1 U5545 ( .B(fifo_array[25]), .A(fifo_array[67]), .S(n5672), .Y(n5099)
         );
  MUX2X1 U5546 ( .B(n5098), .A(n5095), .S(n5727), .Y(n5102) );
  MUX2X1 U5547 ( .B(n5101), .A(n5086), .S(n23), .Y(n5609) );
  MUX2X1 U5548 ( .B(fifo_array[1286]), .A(fifo_array[1328]), .S(n5672), .Y(
        n5106) );
  MUX2X1 U5549 ( .B(fifo_array[1202]), .A(fifo_array[1244]), .S(n5672), .Y(
        n5105) );
  MUX2X1 U5550 ( .B(fifo_array[1118]), .A(fifo_array[1160]), .S(n5672), .Y(
        n5109) );
  MUX2X1 U5551 ( .B(fifo_array[1034]), .A(fifo_array[1076]), .S(n5672), .Y(
        n5108) );
  MUX2X1 U5552 ( .B(n5107), .A(n5104), .S(n5728), .Y(n5118) );
  MUX2X1 U5553 ( .B(fifo_array[950]), .A(fifo_array[992]), .S(n5673), .Y(n5112) );
  MUX2X1 U5554 ( .B(fifo_array[866]), .A(fifo_array[908]), .S(n5673), .Y(n5111) );
  MUX2X1 U5555 ( .B(fifo_array[782]), .A(fifo_array[824]), .S(n5673), .Y(n5115) );
  MUX2X1 U5556 ( .B(fifo_array[698]), .A(fifo_array[740]), .S(n5673), .Y(n5114) );
  MUX2X1 U5557 ( .B(n5113), .A(n5110), .S(n5727), .Y(n5117) );
  MUX2X1 U5558 ( .B(fifo_array[614]), .A(fifo_array[656]), .S(n5673), .Y(n5121) );
  MUX2X1 U5559 ( .B(fifo_array[530]), .A(fifo_array[572]), .S(n5673), .Y(n5120) );
  MUX2X1 U5560 ( .B(fifo_array[446]), .A(fifo_array[488]), .S(n5673), .Y(n5124) );
  MUX2X1 U5561 ( .B(fifo_array[362]), .A(fifo_array[404]), .S(n5673), .Y(n5123) );
  MUX2X1 U5562 ( .B(n5122), .A(n5119), .S(n5729), .Y(n5133) );
  MUX2X1 U5563 ( .B(fifo_array[278]), .A(fifo_array[320]), .S(n5673), .Y(n5127) );
  MUX2X1 U5564 ( .B(fifo_array[194]), .A(fifo_array[236]), .S(n5673), .Y(n5126) );
  MUX2X1 U5565 ( .B(fifo_array[110]), .A(fifo_array[152]), .S(n5673), .Y(n5130) );
  MUX2X1 U5566 ( .B(fifo_array[26]), .A(fifo_array[68]), .S(n5673), .Y(n5129)
         );
  MUX2X1 U5567 ( .B(n5128), .A(n5125), .S(n5726), .Y(n5132) );
  MUX2X1 U5568 ( .B(n5131), .A(n5116), .S(n23), .Y(n5610) );
  MUX2X1 U5569 ( .B(fifo_array[1287]), .A(fifo_array[1329]), .S(n5674), .Y(
        n5136) );
  MUX2X1 U5570 ( .B(fifo_array[1203]), .A(fifo_array[1245]), .S(n5674), .Y(
        n5135) );
  MUX2X1 U5571 ( .B(fifo_array[1119]), .A(fifo_array[1161]), .S(n5674), .Y(
        n5139) );
  MUX2X1 U5572 ( .B(fifo_array[1035]), .A(fifo_array[1077]), .S(n5674), .Y(
        n5138) );
  MUX2X1 U5573 ( .B(n5137), .A(n5134), .S(n21), .Y(n5148) );
  MUX2X1 U5574 ( .B(fifo_array[951]), .A(fifo_array[993]), .S(n5674), .Y(n5142) );
  MUX2X1 U5575 ( .B(fifo_array[867]), .A(fifo_array[909]), .S(n5674), .Y(n5141) );
  MUX2X1 U5576 ( .B(fifo_array[783]), .A(fifo_array[825]), .S(n5674), .Y(n5145) );
  MUX2X1 U5577 ( .B(fifo_array[699]), .A(fifo_array[741]), .S(n5674), .Y(n5144) );
  MUX2X1 U5578 ( .B(n5143), .A(n5140), .S(n21), .Y(n5147) );
  MUX2X1 U5579 ( .B(fifo_array[615]), .A(fifo_array[657]), .S(n5674), .Y(n5151) );
  MUX2X1 U5580 ( .B(fifo_array[531]), .A(fifo_array[573]), .S(n5674), .Y(n5150) );
  MUX2X1 U5581 ( .B(fifo_array[447]), .A(fifo_array[489]), .S(n5674), .Y(n5154) );
  MUX2X1 U5582 ( .B(fifo_array[363]), .A(fifo_array[405]), .S(n5674), .Y(n5153) );
  MUX2X1 U5583 ( .B(n5152), .A(n5149), .S(n21), .Y(n5163) );
  MUX2X1 U5584 ( .B(fifo_array[279]), .A(fifo_array[321]), .S(n5675), .Y(n5157) );
  MUX2X1 U5585 ( .B(fifo_array[195]), .A(fifo_array[237]), .S(n5675), .Y(n5156) );
  MUX2X1 U5586 ( .B(fifo_array[111]), .A(fifo_array[153]), .S(n5675), .Y(n5160) );
  MUX2X1 U5587 ( .B(fifo_array[27]), .A(fifo_array[69]), .S(n5675), .Y(n5159)
         );
  MUX2X1 U5588 ( .B(n5158), .A(n5155), .S(n21), .Y(n5162) );
  MUX2X1 U5589 ( .B(n5161), .A(n5146), .S(n23), .Y(n5611) );
  MUX2X1 U5590 ( .B(fifo_array[1288]), .A(fifo_array[1330]), .S(n5675), .Y(
        n5166) );
  MUX2X1 U5591 ( .B(fifo_array[1204]), .A(fifo_array[1246]), .S(n5675), .Y(
        n5165) );
  MUX2X1 U5592 ( .B(fifo_array[1120]), .A(fifo_array[1162]), .S(n5675), .Y(
        n5169) );
  MUX2X1 U5593 ( .B(fifo_array[1036]), .A(fifo_array[1078]), .S(n5675), .Y(
        n5168) );
  MUX2X1 U5594 ( .B(n5167), .A(n5164), .S(n21), .Y(n5178) );
  MUX2X1 U5595 ( .B(fifo_array[952]), .A(fifo_array[994]), .S(n5675), .Y(n5172) );
  MUX2X1 U5596 ( .B(fifo_array[868]), .A(fifo_array[910]), .S(n5675), .Y(n5171) );
  MUX2X1 U5597 ( .B(fifo_array[784]), .A(fifo_array[826]), .S(n5675), .Y(n5175) );
  MUX2X1 U5598 ( .B(fifo_array[700]), .A(fifo_array[742]), .S(n5675), .Y(n5174) );
  MUX2X1 U5599 ( .B(n5173), .A(n5170), .S(n21), .Y(n5177) );
  MUX2X1 U5600 ( .B(fifo_array[616]), .A(fifo_array[658]), .S(n5676), .Y(n5181) );
  MUX2X1 U5601 ( .B(fifo_array[532]), .A(fifo_array[574]), .S(n5676), .Y(n5180) );
  MUX2X1 U5602 ( .B(fifo_array[448]), .A(fifo_array[490]), .S(n5676), .Y(n5184) );
  MUX2X1 U5603 ( .B(fifo_array[364]), .A(fifo_array[406]), .S(n5676), .Y(n5183) );
  MUX2X1 U5604 ( .B(n5182), .A(n5179), .S(n21), .Y(n5193) );
  MUX2X1 U5605 ( .B(fifo_array[280]), .A(fifo_array[322]), .S(n5676), .Y(n5187) );
  MUX2X1 U5606 ( .B(fifo_array[196]), .A(fifo_array[238]), .S(n5676), .Y(n5186) );
  MUX2X1 U5607 ( .B(fifo_array[112]), .A(fifo_array[154]), .S(n5676), .Y(n5190) );
  MUX2X1 U5608 ( .B(fifo_array[28]), .A(fifo_array[70]), .S(n5676), .Y(n5189)
         );
  MUX2X1 U5609 ( .B(n5188), .A(n5185), .S(n21), .Y(n5192) );
  MUX2X1 U5610 ( .B(n5191), .A(n5176), .S(n23), .Y(n5612) );
  MUX2X1 U5611 ( .B(fifo_array[1289]), .A(fifo_array[1331]), .S(n5676), .Y(
        n5196) );
  MUX2X1 U5612 ( .B(fifo_array[1205]), .A(fifo_array[1247]), .S(n5676), .Y(
        n5195) );
  MUX2X1 U5613 ( .B(fifo_array[1121]), .A(fifo_array[1163]), .S(n5676), .Y(
        n5199) );
  MUX2X1 U5614 ( .B(fifo_array[1037]), .A(fifo_array[1079]), .S(n5676), .Y(
        n5198) );
  MUX2X1 U5615 ( .B(n5197), .A(n5194), .S(n21), .Y(n5208) );
  MUX2X1 U5616 ( .B(fifo_array[953]), .A(fifo_array[995]), .S(n5677), .Y(n5202) );
  MUX2X1 U5617 ( .B(fifo_array[869]), .A(fifo_array[911]), .S(n5677), .Y(n5201) );
  MUX2X1 U5618 ( .B(fifo_array[785]), .A(fifo_array[827]), .S(n5677), .Y(n5205) );
  MUX2X1 U5619 ( .B(fifo_array[701]), .A(fifo_array[743]), .S(n5677), .Y(n5204) );
  MUX2X1 U5620 ( .B(n5203), .A(n5200), .S(n21), .Y(n5207) );
  MUX2X1 U5621 ( .B(fifo_array[617]), .A(fifo_array[659]), .S(n5677), .Y(n5211) );
  MUX2X1 U5622 ( .B(fifo_array[533]), .A(fifo_array[575]), .S(n5677), .Y(n5210) );
  MUX2X1 U5623 ( .B(fifo_array[449]), .A(fifo_array[491]), .S(n5677), .Y(n5214) );
  MUX2X1 U5624 ( .B(fifo_array[365]), .A(fifo_array[407]), .S(n5677), .Y(n5213) );
  MUX2X1 U5625 ( .B(n5212), .A(n5209), .S(n21), .Y(n5223) );
  MUX2X1 U5626 ( .B(fifo_array[281]), .A(fifo_array[323]), .S(n5677), .Y(n5217) );
  MUX2X1 U5627 ( .B(fifo_array[197]), .A(fifo_array[239]), .S(n5677), .Y(n5216) );
  MUX2X1 U5628 ( .B(fifo_array[113]), .A(fifo_array[155]), .S(n5677), .Y(n5220) );
  MUX2X1 U5629 ( .B(fifo_array[29]), .A(fifo_array[71]), .S(n5677), .Y(n5219)
         );
  MUX2X1 U5630 ( .B(n5218), .A(n5215), .S(n21), .Y(n5222) );
  MUX2X1 U5631 ( .B(n5221), .A(n5206), .S(n23), .Y(n5613) );
  MUX2X1 U5632 ( .B(fifo_array[1290]), .A(fifo_array[1332]), .S(n5678), .Y(
        n5226) );
  MUX2X1 U5633 ( .B(fifo_array[1206]), .A(fifo_array[1248]), .S(n5678), .Y(
        n5225) );
  MUX2X1 U5634 ( .B(fifo_array[1122]), .A(fifo_array[1164]), .S(n5678), .Y(
        n5229) );
  MUX2X1 U5635 ( .B(fifo_array[1038]), .A(fifo_array[1080]), .S(n5678), .Y(
        n5228) );
  MUX2X1 U5636 ( .B(n5227), .A(n5224), .S(n21), .Y(n5238) );
  MUX2X1 U5637 ( .B(fifo_array[954]), .A(fifo_array[996]), .S(n5678), .Y(n5232) );
  MUX2X1 U5638 ( .B(fifo_array[870]), .A(fifo_array[912]), .S(n5678), .Y(n5231) );
  MUX2X1 U5639 ( .B(fifo_array[786]), .A(fifo_array[828]), .S(n5678), .Y(n5235) );
  MUX2X1 U5640 ( .B(fifo_array[702]), .A(fifo_array[744]), .S(n5678), .Y(n5234) );
  MUX2X1 U5641 ( .B(n5233), .A(n5230), .S(n21), .Y(n5237) );
  MUX2X1 U5642 ( .B(fifo_array[618]), .A(fifo_array[660]), .S(n5678), .Y(n5241) );
  MUX2X1 U5643 ( .B(fifo_array[534]), .A(fifo_array[576]), .S(n5678), .Y(n5240) );
  MUX2X1 U5644 ( .B(fifo_array[450]), .A(fifo_array[492]), .S(n5678), .Y(n5244) );
  MUX2X1 U5645 ( .B(fifo_array[366]), .A(fifo_array[408]), .S(n5678), .Y(n5243) );
  MUX2X1 U5646 ( .B(n5242), .A(n5239), .S(n21), .Y(n5253) );
  MUX2X1 U5647 ( .B(fifo_array[282]), .A(fifo_array[324]), .S(n5679), .Y(n5247) );
  MUX2X1 U5648 ( .B(fifo_array[198]), .A(fifo_array[240]), .S(n5679), .Y(n5246) );
  MUX2X1 U5649 ( .B(fifo_array[114]), .A(fifo_array[156]), .S(n5679), .Y(n5250) );
  MUX2X1 U5650 ( .B(fifo_array[30]), .A(fifo_array[72]), .S(n5679), .Y(n5249)
         );
  MUX2X1 U5651 ( .B(n5248), .A(n5245), .S(n21), .Y(n5252) );
  MUX2X1 U5652 ( .B(n5251), .A(n5236), .S(n23), .Y(n5614) );
  MUX2X1 U5653 ( .B(fifo_array[1291]), .A(fifo_array[1333]), .S(n5679), .Y(
        n5256) );
  MUX2X1 U5654 ( .B(fifo_array[1207]), .A(fifo_array[1249]), .S(n5679), .Y(
        n5255) );
  MUX2X1 U5655 ( .B(fifo_array[1123]), .A(fifo_array[1165]), .S(n5679), .Y(
        n5259) );
  MUX2X1 U5656 ( .B(fifo_array[1039]), .A(fifo_array[1081]), .S(n5679), .Y(
        n5258) );
  MUX2X1 U5657 ( .B(n5257), .A(n5254), .S(n21), .Y(n5268) );
  MUX2X1 U5658 ( .B(fifo_array[955]), .A(fifo_array[997]), .S(n5679), .Y(n5262) );
  MUX2X1 U5659 ( .B(fifo_array[871]), .A(fifo_array[913]), .S(n5679), .Y(n5261) );
  MUX2X1 U5660 ( .B(fifo_array[787]), .A(fifo_array[829]), .S(n5679), .Y(n5265) );
  MUX2X1 U5661 ( .B(fifo_array[703]), .A(fifo_array[745]), .S(n5679), .Y(n5264) );
  MUX2X1 U5662 ( .B(n5263), .A(n5260), .S(n21), .Y(n5267) );
  MUX2X1 U5663 ( .B(fifo_array[619]), .A(fifo_array[661]), .S(n5680), .Y(n5271) );
  MUX2X1 U5664 ( .B(fifo_array[535]), .A(fifo_array[577]), .S(n5680), .Y(n5270) );
  MUX2X1 U5665 ( .B(fifo_array[451]), .A(fifo_array[493]), .S(n5680), .Y(n5274) );
  MUX2X1 U5666 ( .B(fifo_array[367]), .A(fifo_array[409]), .S(n5680), .Y(n5273) );
  MUX2X1 U5667 ( .B(n5272), .A(n5269), .S(n21), .Y(n5283) );
  MUX2X1 U5668 ( .B(fifo_array[283]), .A(fifo_array[325]), .S(n5680), .Y(n5277) );
  MUX2X1 U5669 ( .B(fifo_array[199]), .A(fifo_array[241]), .S(n5680), .Y(n5276) );
  MUX2X1 U5670 ( .B(fifo_array[115]), .A(fifo_array[157]), .S(n5680), .Y(n5280) );
  MUX2X1 U5671 ( .B(fifo_array[31]), .A(fifo_array[73]), .S(n5680), .Y(n5279)
         );
  MUX2X1 U5672 ( .B(n5278), .A(n5275), .S(n21), .Y(n5282) );
  MUX2X1 U5673 ( .B(n5281), .A(n5266), .S(n23), .Y(n5615) );
  MUX2X1 U5674 ( .B(fifo_array[1292]), .A(fifo_array[1334]), .S(n5680), .Y(
        n5286) );
  MUX2X1 U5675 ( .B(fifo_array[1208]), .A(fifo_array[1250]), .S(n5680), .Y(
        n5285) );
  MUX2X1 U5676 ( .B(fifo_array[1124]), .A(fifo_array[1166]), .S(n5680), .Y(
        n5289) );
  MUX2X1 U5677 ( .B(fifo_array[1040]), .A(fifo_array[1082]), .S(n5680), .Y(
        n5288) );
  MUX2X1 U5678 ( .B(n5287), .A(n5284), .S(n21), .Y(n5298) );
  MUX2X1 U5679 ( .B(fifo_array[956]), .A(fifo_array[998]), .S(n5681), .Y(n5292) );
  MUX2X1 U5680 ( .B(fifo_array[872]), .A(fifo_array[914]), .S(n5681), .Y(n5291) );
  MUX2X1 U5681 ( .B(fifo_array[788]), .A(fifo_array[830]), .S(n5681), .Y(n5295) );
  MUX2X1 U5682 ( .B(fifo_array[704]), .A(fifo_array[746]), .S(n5681), .Y(n5294) );
  MUX2X1 U5683 ( .B(n5293), .A(n5290), .S(n21), .Y(n5297) );
  MUX2X1 U5684 ( .B(fifo_array[620]), .A(fifo_array[662]), .S(n5681), .Y(n5301) );
  MUX2X1 U5685 ( .B(fifo_array[536]), .A(fifo_array[578]), .S(n5681), .Y(n5300) );
  MUX2X1 U5686 ( .B(fifo_array[452]), .A(fifo_array[494]), .S(n5681), .Y(n5304) );
  MUX2X1 U5687 ( .B(fifo_array[368]), .A(fifo_array[410]), .S(n5681), .Y(n5303) );
  MUX2X1 U5688 ( .B(n5302), .A(n5299), .S(n21), .Y(n5313) );
  MUX2X1 U5689 ( .B(fifo_array[284]), .A(fifo_array[326]), .S(n5681), .Y(n5307) );
  MUX2X1 U5690 ( .B(fifo_array[200]), .A(fifo_array[242]), .S(n5681), .Y(n5306) );
  MUX2X1 U5691 ( .B(fifo_array[116]), .A(fifo_array[158]), .S(n5681), .Y(n5310) );
  MUX2X1 U5692 ( .B(fifo_array[32]), .A(fifo_array[74]), .S(n5681), .Y(n5309)
         );
  MUX2X1 U5693 ( .B(n5308), .A(n5305), .S(n21), .Y(n5312) );
  MUX2X1 U5694 ( .B(n5311), .A(n5296), .S(n23), .Y(n5616) );
  MUX2X1 U5695 ( .B(fifo_array[1293]), .A(fifo_array[1335]), .S(n5682), .Y(
        n5316) );
  MUX2X1 U5696 ( .B(fifo_array[1209]), .A(fifo_array[1251]), .S(n5682), .Y(
        n5315) );
  MUX2X1 U5697 ( .B(fifo_array[1125]), .A(fifo_array[1167]), .S(n5682), .Y(
        n5319) );
  MUX2X1 U5698 ( .B(fifo_array[1041]), .A(fifo_array[1083]), .S(n5682), .Y(
        n5318) );
  MUX2X1 U5699 ( .B(n5317), .A(n5314), .S(n5730), .Y(n5328) );
  MUX2X1 U5700 ( .B(fifo_array[957]), .A(fifo_array[999]), .S(n5682), .Y(n5322) );
  MUX2X1 U5701 ( .B(fifo_array[873]), .A(fifo_array[915]), .S(n5682), .Y(n5321) );
  MUX2X1 U5702 ( .B(fifo_array[789]), .A(fifo_array[831]), .S(n5682), .Y(n5325) );
  MUX2X1 U5703 ( .B(fifo_array[705]), .A(fifo_array[747]), .S(n5682), .Y(n5324) );
  MUX2X1 U5704 ( .B(n5323), .A(n5320), .S(n21), .Y(n5327) );
  MUX2X1 U5705 ( .B(fifo_array[621]), .A(fifo_array[663]), .S(n5682), .Y(n5331) );
  MUX2X1 U5706 ( .B(fifo_array[537]), .A(fifo_array[579]), .S(n5682), .Y(n5330) );
  MUX2X1 U5707 ( .B(fifo_array[453]), .A(fifo_array[495]), .S(n5682), .Y(n5334) );
  MUX2X1 U5708 ( .B(fifo_array[369]), .A(fifo_array[411]), .S(n5682), .Y(n5333) );
  MUX2X1 U5709 ( .B(n5332), .A(n5329), .S(n21), .Y(n5343) );
  MUX2X1 U5710 ( .B(fifo_array[285]), .A(fifo_array[327]), .S(n5683), .Y(n5337) );
  MUX2X1 U5711 ( .B(fifo_array[201]), .A(fifo_array[243]), .S(n5683), .Y(n5336) );
  MUX2X1 U5712 ( .B(fifo_array[117]), .A(fifo_array[159]), .S(n5683), .Y(n5340) );
  MUX2X1 U5713 ( .B(fifo_array[33]), .A(fifo_array[75]), .S(n5683), .Y(n5339)
         );
  MUX2X1 U5714 ( .B(n5338), .A(n5335), .S(n21), .Y(n5342) );
  MUX2X1 U5715 ( .B(n5341), .A(n5326), .S(n23), .Y(n5617) );
  MUX2X1 U5716 ( .B(fifo_array[1294]), .A(fifo_array[1336]), .S(n5683), .Y(
        n5346) );
  MUX2X1 U5717 ( .B(fifo_array[1210]), .A(fifo_array[1252]), .S(n5683), .Y(
        n5345) );
  MUX2X1 U5718 ( .B(fifo_array[1126]), .A(fifo_array[1168]), .S(n5683), .Y(
        n5349) );
  MUX2X1 U5719 ( .B(fifo_array[1042]), .A(fifo_array[1084]), .S(n5683), .Y(
        n5348) );
  MUX2X1 U5720 ( .B(n5347), .A(n5344), .S(n21), .Y(n5358) );
  MUX2X1 U5721 ( .B(fifo_array[958]), .A(fifo_array[1000]), .S(n5683), .Y(
        n5352) );
  MUX2X1 U5722 ( .B(fifo_array[874]), .A(fifo_array[916]), .S(n5683), .Y(n5351) );
  MUX2X1 U5723 ( .B(fifo_array[790]), .A(fifo_array[832]), .S(n5683), .Y(n5355) );
  MUX2X1 U5724 ( .B(fifo_array[706]), .A(fifo_array[748]), .S(n5683), .Y(n5354) );
  MUX2X1 U5725 ( .B(n5353), .A(n5350), .S(n5730), .Y(n5357) );
  MUX2X1 U5726 ( .B(fifo_array[622]), .A(fifo_array[664]), .S(n5684), .Y(n5361) );
  MUX2X1 U5727 ( .B(fifo_array[538]), .A(fifo_array[580]), .S(n5684), .Y(n5360) );
  MUX2X1 U5728 ( .B(fifo_array[454]), .A(fifo_array[496]), .S(n5684), .Y(n5364) );
  MUX2X1 U5729 ( .B(fifo_array[370]), .A(fifo_array[412]), .S(n5684), .Y(n5363) );
  MUX2X1 U5730 ( .B(n5362), .A(n5359), .S(n21), .Y(n5373) );
  MUX2X1 U5731 ( .B(fifo_array[286]), .A(fifo_array[328]), .S(n5684), .Y(n5367) );
  MUX2X1 U5732 ( .B(fifo_array[202]), .A(fifo_array[244]), .S(n5684), .Y(n5366) );
  MUX2X1 U5733 ( .B(fifo_array[118]), .A(fifo_array[160]), .S(n5684), .Y(n5370) );
  MUX2X1 U5734 ( .B(fifo_array[34]), .A(fifo_array[76]), .S(n5684), .Y(n5369)
         );
  MUX2X1 U5735 ( .B(n5368), .A(n5365), .S(n21), .Y(n5372) );
  MUX2X1 U5736 ( .B(n5371), .A(n5356), .S(n23), .Y(n5618) );
  MUX2X1 U5737 ( .B(fifo_array[1295]), .A(fifo_array[1337]), .S(n5684), .Y(
        n5376) );
  MUX2X1 U5738 ( .B(fifo_array[1211]), .A(fifo_array[1253]), .S(n5684), .Y(
        n5375) );
  MUX2X1 U5739 ( .B(fifo_array[1127]), .A(fifo_array[1169]), .S(n5684), .Y(
        n5379) );
  MUX2X1 U5740 ( .B(fifo_array[1043]), .A(fifo_array[1085]), .S(n5684), .Y(
        n5378) );
  MUX2X1 U5741 ( .B(n5377), .A(n5374), .S(n21), .Y(n5388) );
  MUX2X1 U5742 ( .B(fifo_array[959]), .A(fifo_array[1001]), .S(n5685), .Y(
        n5382) );
  MUX2X1 U5743 ( .B(fifo_array[875]), .A(fifo_array[917]), .S(n5685), .Y(n5381) );
  MUX2X1 U5744 ( .B(fifo_array[791]), .A(fifo_array[833]), .S(n5685), .Y(n5385) );
  MUX2X1 U5745 ( .B(fifo_array[707]), .A(fifo_array[749]), .S(n5685), .Y(n5384) );
  MUX2X1 U5746 ( .B(n5383), .A(n5380), .S(n21), .Y(n5387) );
  MUX2X1 U5747 ( .B(fifo_array[623]), .A(fifo_array[665]), .S(n5685), .Y(n5391) );
  MUX2X1 U5748 ( .B(fifo_array[539]), .A(fifo_array[581]), .S(n5685), .Y(n5390) );
  MUX2X1 U5749 ( .B(fifo_array[455]), .A(fifo_array[497]), .S(n5685), .Y(n5394) );
  MUX2X1 U5750 ( .B(fifo_array[371]), .A(fifo_array[413]), .S(n5685), .Y(n5393) );
  MUX2X1 U5751 ( .B(n5392), .A(n5389), .S(n5730), .Y(n5403) );
  MUX2X1 U5752 ( .B(fifo_array[287]), .A(fifo_array[329]), .S(n5685), .Y(n5397) );
  MUX2X1 U5753 ( .B(fifo_array[203]), .A(fifo_array[245]), .S(n5685), .Y(n5396) );
  MUX2X1 U5754 ( .B(fifo_array[119]), .A(fifo_array[161]), .S(n5685), .Y(n5400) );
  MUX2X1 U5755 ( .B(fifo_array[35]), .A(fifo_array[77]), .S(n5685), .Y(n5399)
         );
  MUX2X1 U5756 ( .B(n5398), .A(n5395), .S(n21), .Y(n5402) );
  MUX2X1 U5757 ( .B(n5401), .A(n5386), .S(n23), .Y(n5619) );
  MUX2X1 U5758 ( .B(fifo_array[1296]), .A(fifo_array[1338]), .S(n5686), .Y(
        n5406) );
  MUX2X1 U5759 ( .B(fifo_array[1212]), .A(fifo_array[1254]), .S(n5686), .Y(
        n5405) );
  MUX2X1 U5760 ( .B(fifo_array[1128]), .A(fifo_array[1170]), .S(n5686), .Y(
        n5409) );
  MUX2X1 U5761 ( .B(fifo_array[1044]), .A(fifo_array[1086]), .S(n5686), .Y(
        n5408) );
  MUX2X1 U5762 ( .B(n5407), .A(n5404), .S(n21), .Y(n5418) );
  MUX2X1 U5763 ( .B(fifo_array[960]), .A(fifo_array[1002]), .S(n5686), .Y(
        n5412) );
  MUX2X1 U5764 ( .B(fifo_array[876]), .A(fifo_array[918]), .S(n5686), .Y(n5411) );
  MUX2X1 U5765 ( .B(fifo_array[792]), .A(fifo_array[834]), .S(n5686), .Y(n5415) );
  MUX2X1 U5766 ( .B(fifo_array[708]), .A(fifo_array[750]), .S(n5686), .Y(n5414) );
  MUX2X1 U5767 ( .B(n5413), .A(n5410), .S(n21), .Y(n5417) );
  MUX2X1 U5768 ( .B(fifo_array[624]), .A(fifo_array[666]), .S(n5686), .Y(n5421) );
  MUX2X1 U5769 ( .B(fifo_array[540]), .A(fifo_array[582]), .S(n5686), .Y(n5420) );
  MUX2X1 U5770 ( .B(fifo_array[456]), .A(fifo_array[498]), .S(n5686), .Y(n5424) );
  MUX2X1 U5771 ( .B(fifo_array[372]), .A(fifo_array[414]), .S(n5686), .Y(n5423) );
  MUX2X1 U5772 ( .B(n5422), .A(n5419), .S(n21), .Y(n5433) );
  MUX2X1 U5773 ( .B(fifo_array[288]), .A(fifo_array[330]), .S(n5687), .Y(n5427) );
  MUX2X1 U5774 ( .B(fifo_array[204]), .A(fifo_array[246]), .S(n5687), .Y(n5426) );
  MUX2X1 U5775 ( .B(fifo_array[120]), .A(fifo_array[162]), .S(n5687), .Y(n5430) );
  MUX2X1 U5776 ( .B(fifo_array[36]), .A(fifo_array[78]), .S(n5687), .Y(n5429)
         );
  MUX2X1 U5777 ( .B(n5428), .A(n5425), .S(n21), .Y(n5432) );
  MUX2X1 U5778 ( .B(n5431), .A(n5416), .S(n23), .Y(n5620) );
  MUX2X1 U5779 ( .B(fifo_array[1297]), .A(fifo_array[1339]), .S(n5687), .Y(
        n5436) );
  MUX2X1 U5780 ( .B(fifo_array[1213]), .A(fifo_array[1255]), .S(n5687), .Y(
        n5435) );
  MUX2X1 U5781 ( .B(fifo_array[1129]), .A(fifo_array[1171]), .S(n5687), .Y(
        n5439) );
  MUX2X1 U5782 ( .B(fifo_array[1045]), .A(fifo_array[1087]), .S(n5687), .Y(
        n5438) );
  MUX2X1 U5783 ( .B(n5437), .A(n5434), .S(n21), .Y(n5448) );
  MUX2X1 U5784 ( .B(fifo_array[961]), .A(fifo_array[1003]), .S(n5687), .Y(
        n5442) );
  MUX2X1 U5785 ( .B(fifo_array[877]), .A(fifo_array[919]), .S(n5687), .Y(n5441) );
  MUX2X1 U5786 ( .B(fifo_array[793]), .A(fifo_array[835]), .S(n5687), .Y(n5445) );
  MUX2X1 U5787 ( .B(fifo_array[709]), .A(fifo_array[751]), .S(n5687), .Y(n5444) );
  MUX2X1 U5788 ( .B(n5443), .A(n5440), .S(n21), .Y(n5447) );
  MUX2X1 U5789 ( .B(fifo_array[625]), .A(fifo_array[667]), .S(n5688), .Y(n5451) );
  MUX2X1 U5790 ( .B(fifo_array[541]), .A(fifo_array[583]), .S(n5688), .Y(n5450) );
  MUX2X1 U5791 ( .B(fifo_array[457]), .A(fifo_array[499]), .S(n5688), .Y(n5454) );
  MUX2X1 U5792 ( .B(fifo_array[373]), .A(fifo_array[415]), .S(n5688), .Y(n5453) );
  MUX2X1 U5793 ( .B(n5452), .A(n5449), .S(n21), .Y(n5463) );
  MUX2X1 U5794 ( .B(fifo_array[289]), .A(fifo_array[331]), .S(n5688), .Y(n5457) );
  MUX2X1 U5795 ( .B(fifo_array[205]), .A(fifo_array[247]), .S(n5688), .Y(n5456) );
  MUX2X1 U5796 ( .B(fifo_array[121]), .A(fifo_array[163]), .S(n5688), .Y(n5460) );
  MUX2X1 U5797 ( .B(fifo_array[37]), .A(fifo_array[79]), .S(n5688), .Y(n5459)
         );
  MUX2X1 U5798 ( .B(n5458), .A(n5455), .S(n21), .Y(n5462) );
  MUX2X1 U5799 ( .B(n5461), .A(n5446), .S(n23), .Y(n5621) );
  MUX2X1 U5800 ( .B(fifo_array[1298]), .A(fifo_array[1340]), .S(n5688), .Y(
        n5466) );
  MUX2X1 U5801 ( .B(fifo_array[1214]), .A(fifo_array[1256]), .S(n5688), .Y(
        n5465) );
  MUX2X1 U5802 ( .B(fifo_array[1130]), .A(fifo_array[1172]), .S(n5688), .Y(
        n5469) );
  MUX2X1 U5803 ( .B(fifo_array[1046]), .A(fifo_array[1088]), .S(n5688), .Y(
        n5468) );
  MUX2X1 U5804 ( .B(n5467), .A(n5464), .S(n21), .Y(n5478) );
  MUX2X1 U5805 ( .B(fifo_array[962]), .A(fifo_array[1004]), .S(n5689), .Y(
        n5472) );
  MUX2X1 U5806 ( .B(fifo_array[878]), .A(fifo_array[920]), .S(n5689), .Y(n5471) );
  MUX2X1 U5807 ( .B(fifo_array[794]), .A(fifo_array[836]), .S(n5689), .Y(n5475) );
  MUX2X1 U5808 ( .B(fifo_array[710]), .A(fifo_array[752]), .S(n5689), .Y(n5474) );
  MUX2X1 U5809 ( .B(n5473), .A(n5470), .S(n21), .Y(n5477) );
  MUX2X1 U5810 ( .B(fifo_array[626]), .A(fifo_array[668]), .S(n5689), .Y(n5481) );
  MUX2X1 U5811 ( .B(fifo_array[542]), .A(fifo_array[584]), .S(n5689), .Y(n5480) );
  MUX2X1 U5812 ( .B(fifo_array[458]), .A(fifo_array[500]), .S(n5689), .Y(n5484) );
  MUX2X1 U5813 ( .B(fifo_array[374]), .A(fifo_array[416]), .S(n5689), .Y(n5483) );
  MUX2X1 U5814 ( .B(n5482), .A(n5479), .S(n21), .Y(n5493) );
  MUX2X1 U5815 ( .B(fifo_array[290]), .A(fifo_array[332]), .S(n5689), .Y(n5487) );
  MUX2X1 U5816 ( .B(fifo_array[206]), .A(fifo_array[248]), .S(n5689), .Y(n5486) );
  MUX2X1 U5817 ( .B(fifo_array[122]), .A(fifo_array[164]), .S(n5689), .Y(n5490) );
  MUX2X1 U5818 ( .B(fifo_array[38]), .A(fifo_array[80]), .S(n5689), .Y(n5489)
         );
  MUX2X1 U5819 ( .B(n5488), .A(n5485), .S(n21), .Y(n5492) );
  MUX2X1 U5820 ( .B(n5491), .A(n5476), .S(n23), .Y(n5622) );
  MUX2X1 U5821 ( .B(fifo_array[1299]), .A(fifo_array[1341]), .S(n5690), .Y(
        n5496) );
  MUX2X1 U5822 ( .B(fifo_array[1215]), .A(fifo_array[1257]), .S(n5690), .Y(
        n5495) );
  MUX2X1 U5823 ( .B(fifo_array[1131]), .A(fifo_array[1173]), .S(n5690), .Y(
        n5499) );
  MUX2X1 U5824 ( .B(fifo_array[1047]), .A(fifo_array[1089]), .S(n5690), .Y(
        n5498) );
  MUX2X1 U5825 ( .B(n5497), .A(n5494), .S(n5730), .Y(n5508) );
  MUX2X1 U5826 ( .B(fifo_array[963]), .A(fifo_array[1005]), .S(n5690), .Y(
        n5502) );
  MUX2X1 U5827 ( .B(fifo_array[879]), .A(fifo_array[921]), .S(n5690), .Y(n5501) );
  MUX2X1 U5828 ( .B(fifo_array[795]), .A(fifo_array[837]), .S(n5690), .Y(n5505) );
  MUX2X1 U5829 ( .B(fifo_array[711]), .A(fifo_array[753]), .S(n5690), .Y(n5504) );
  MUX2X1 U5830 ( .B(n5503), .A(n5500), .S(n5730), .Y(n5507) );
  MUX2X1 U5831 ( .B(fifo_array[627]), .A(fifo_array[669]), .S(n5690), .Y(n5511) );
  MUX2X1 U5832 ( .B(fifo_array[543]), .A(fifo_array[585]), .S(n5690), .Y(n5510) );
  MUX2X1 U5833 ( .B(fifo_array[459]), .A(fifo_array[501]), .S(n5690), .Y(n5514) );
  MUX2X1 U5834 ( .B(fifo_array[375]), .A(fifo_array[417]), .S(n5690), .Y(n5513) );
  MUX2X1 U5835 ( .B(n5512), .A(n5509), .S(n5730), .Y(n5523) );
  MUX2X1 U5836 ( .B(fifo_array[291]), .A(fifo_array[333]), .S(n5691), .Y(n5517) );
  MUX2X1 U5837 ( .B(fifo_array[207]), .A(fifo_array[249]), .S(n5691), .Y(n5516) );
  MUX2X1 U5838 ( .B(fifo_array[123]), .A(fifo_array[165]), .S(n5691), .Y(n5520) );
  MUX2X1 U5839 ( .B(fifo_array[39]), .A(fifo_array[81]), .S(n5691), .Y(n5519)
         );
  MUX2X1 U5840 ( .B(n5518), .A(n5515), .S(n5730), .Y(n5522) );
  MUX2X1 U5841 ( .B(n5521), .A(n5506), .S(n23), .Y(n5623) );
  MUX2X1 U5842 ( .B(fifo_array[1300]), .A(fifo_array[1342]), .S(n5691), .Y(
        n5526) );
  MUX2X1 U5843 ( .B(fifo_array[1216]), .A(fifo_array[1258]), .S(n5691), .Y(
        n5525) );
  MUX2X1 U5844 ( .B(fifo_array[1132]), .A(fifo_array[1174]), .S(n5691), .Y(
        n5529) );
  MUX2X1 U5845 ( .B(fifo_array[1048]), .A(fifo_array[1090]), .S(n5691), .Y(
        n5528) );
  MUX2X1 U5846 ( .B(n5527), .A(n5524), .S(n5730), .Y(n5538) );
  MUX2X1 U5847 ( .B(fifo_array[964]), .A(fifo_array[1006]), .S(n5691), .Y(
        n5532) );
  MUX2X1 U5848 ( .B(fifo_array[880]), .A(fifo_array[922]), .S(n5691), .Y(n5531) );
  MUX2X1 U5849 ( .B(fifo_array[796]), .A(fifo_array[838]), .S(n5691), .Y(n5535) );
  MUX2X1 U5850 ( .B(fifo_array[712]), .A(fifo_array[754]), .S(n5691), .Y(n5534) );
  MUX2X1 U5851 ( .B(n5533), .A(n5530), .S(n5730), .Y(n5537) );
  MUX2X1 U5852 ( .B(fifo_array[628]), .A(fifo_array[670]), .S(n5692), .Y(n5541) );
  MUX2X1 U5853 ( .B(fifo_array[544]), .A(fifo_array[586]), .S(n5692), .Y(n5540) );
  MUX2X1 U5854 ( .B(fifo_array[460]), .A(fifo_array[502]), .S(n5692), .Y(n5544) );
  MUX2X1 U5855 ( .B(fifo_array[376]), .A(fifo_array[418]), .S(n5692), .Y(n5543) );
  MUX2X1 U5856 ( .B(n5542), .A(n5539), .S(n5730), .Y(n5553) );
  MUX2X1 U5857 ( .B(fifo_array[292]), .A(fifo_array[334]), .S(n5692), .Y(n5547) );
  MUX2X1 U5858 ( .B(fifo_array[208]), .A(fifo_array[250]), .S(n5692), .Y(n5546) );
  MUX2X1 U5859 ( .B(fifo_array[124]), .A(fifo_array[166]), .S(n5692), .Y(n5550) );
  MUX2X1 U5860 ( .B(fifo_array[40]), .A(fifo_array[82]), .S(n5692), .Y(n5549)
         );
  MUX2X1 U5861 ( .B(n5548), .A(n5545), .S(n5730), .Y(n5552) );
  MUX2X1 U5862 ( .B(n5551), .A(n5536), .S(n23), .Y(n5624) );
  MUX2X1 U5863 ( .B(fifo_array[1301]), .A(fifo_array[1343]), .S(n5692), .Y(
        n5556) );
  MUX2X1 U5864 ( .B(fifo_array[1217]), .A(fifo_array[1259]), .S(n5692), .Y(
        n5555) );
  MUX2X1 U5865 ( .B(fifo_array[1133]), .A(fifo_array[1175]), .S(n5692), .Y(
        n5559) );
  MUX2X1 U5866 ( .B(fifo_array[1049]), .A(fifo_array[1091]), .S(n5692), .Y(
        n5558) );
  MUX2X1 U5867 ( .B(n5557), .A(n5554), .S(n5730), .Y(n5568) );
  MUX2X1 U5868 ( .B(fifo_array[965]), .A(fifo_array[1007]), .S(n5693), .Y(
        n5562) );
  MUX2X1 U5869 ( .B(fifo_array[881]), .A(fifo_array[923]), .S(n5693), .Y(n5561) );
  MUX2X1 U5870 ( .B(fifo_array[797]), .A(fifo_array[839]), .S(n5693), .Y(n5565) );
  MUX2X1 U5871 ( .B(fifo_array[713]), .A(fifo_array[755]), .S(n5693), .Y(n5564) );
  MUX2X1 U5872 ( .B(n5563), .A(n5560), .S(n5730), .Y(n5567) );
  MUX2X1 U5873 ( .B(fifo_array[629]), .A(fifo_array[671]), .S(n5693), .Y(n5571) );
  MUX2X1 U5874 ( .B(fifo_array[545]), .A(fifo_array[587]), .S(n5693), .Y(n5570) );
  MUX2X1 U5875 ( .B(fifo_array[461]), .A(fifo_array[503]), .S(n5693), .Y(n5574) );
  MUX2X1 U5876 ( .B(fifo_array[377]), .A(fifo_array[419]), .S(n5693), .Y(n5573) );
  MUX2X1 U5877 ( .B(n5572), .A(n5569), .S(n5730), .Y(n5583) );
  MUX2X1 U5878 ( .B(fifo_array[293]), .A(fifo_array[335]), .S(n5693), .Y(n5577) );
  MUX2X1 U5879 ( .B(fifo_array[209]), .A(fifo_array[251]), .S(n5693), .Y(n5576) );
  MUX2X1 U5880 ( .B(fifo_array[125]), .A(fifo_array[167]), .S(n5693), .Y(n5580) );
  MUX2X1 U5881 ( .B(fifo_array[41]), .A(fifo_array[83]), .S(n5693), .Y(n5579)
         );
  MUX2X1 U5882 ( .B(n5578), .A(n5575), .S(n5730), .Y(n5582) );
  MUX2X1 U5883 ( .B(n5581), .A(n5566), .S(n23), .Y(n5625) );
  XOR2X1 U5884 ( .A(r307_carry[4]), .B(wr_ptr[4]), .Y(n79) );
  XOR2X1 U5885 ( .A(r308_carry[4]), .B(n23), .Y(n84) );
  XOR2X1 U5886 ( .A(add_45_carry[5]), .B(fillcount[5]), .Y(n96) );
  OAI21X1 U5887 ( .A(n103), .B(n5904), .C(n4319), .Y(n104) );
  OAI21X1 U5888 ( .A(n5846), .B(n5851), .C(n4229), .Y(n105) );
  OAI21X1 U5889 ( .A(n5847), .B(n5850), .C(n4320), .Y(n106) );
  XNOR2X1 U5890 ( .A(fillcount[4]), .B(n4320), .Y(n107) );
  XNOR2X1 U5891 ( .A(fillcount[5]), .B(n5849), .Y(n108) );
endmodule


module ddr3_init_engine_DW01_inc_0 ( A, SUM );
  input [18:0] A;
  output [18:0] SUM;

  wire   [18:2] carry;

  HAX1 U1_1_17 ( .A(A[17]), .B(carry[17]), .YC(carry[18]), .YS(SUM[17]) );
  HAX1 U1_1_16 ( .A(A[16]), .B(carry[16]), .YC(carry[17]), .YS(SUM[16]) );
  HAX1 U1_1_15 ( .A(A[15]), .B(carry[15]), .YC(carry[16]), .YS(SUM[15]) );
  HAX1 U1_1_14 ( .A(A[14]), .B(carry[14]), .YC(carry[15]), .YS(SUM[14]) );
  HAX1 U1_1_13 ( .A(A[13]), .B(carry[13]), .YC(carry[14]), .YS(SUM[13]) );
  HAX1 U1_1_12 ( .A(A[12]), .B(carry[12]), .YC(carry[13]), .YS(SUM[12]) );
  HAX1 U1_1_11 ( .A(A[11]), .B(carry[11]), .YC(carry[12]), .YS(SUM[11]) );
  HAX1 U1_1_10 ( .A(A[10]), .B(carry[10]), .YC(carry[11]), .YS(SUM[10]) );
  HAX1 U1_1_9 ( .A(A[9]), .B(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  HAX1 U1_1_8 ( .A(A[8]), .B(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  HAX1 U1_1_7 ( .A(A[7]), .B(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[18]), .B(A[18]), .Y(SUM[18]) );
endmodule


module ddr3_init_engine ( ready, csbar, rasbar, casbar, webar, ba, a, odt, 
        ts_con, cke, resetbar, clk, reset, init, ck );
  output [2:0] ba;
  output [12:0] a;
  input clk, reset, init, ck;
  output ready, csbar, rasbar, casbar, webar, odt, ts_con, cke, resetbar;
  wire   flag, RESET, INIT, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n346, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n1, n2,
         n3, n4, n5, n6, n7, n8, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n143, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286;
  wire   [18:0] counter;
  assign csbar = 1'b0;
  assign ba[2] = 1'b0;
  assign a[12] = 1'b0;
  assign a[11] = 1'b0;
  assign a[9] = 1'b0;
  assign a[7] = 1'b0;
  assign a[6] = 1'b0;
  assign a[5] = 1'b0;
  assign a[3] = 1'b0;
  assign a[2] = 1'b0;
  assign a[1] = 1'b0;
  assign a[0] = 1'b0;
  assign odt = 1'b0;
  assign ts_con = 1'b0;

  DFFPOSX1 RESET_reg ( .D(reset), .CLK(clk), .Q(RESET) );
  DFFPOSX1 INIT_reg ( .D(init), .CLK(clk), .Q(INIT) );
  DFFPOSX1 flag_reg ( .D(n249), .CLK(clk), .Q(flag) );
  DFFPOSX1 counter_reg_0_ ( .D(n190), .CLK(clk), .Q(counter[0]) );
  DFFPOSX1 counter_reg_1_ ( .D(n189), .CLK(clk), .Q(counter[1]) );
  DFFPOSX1 counter_reg_2_ ( .D(n188), .CLK(clk), .Q(counter[2]) );
  DFFPOSX1 counter_reg_3_ ( .D(n187), .CLK(clk), .Q(counter[3]) );
  DFFPOSX1 counter_reg_4_ ( .D(n186), .CLK(clk), .Q(counter[4]) );
  DFFPOSX1 counter_reg_5_ ( .D(n185), .CLK(clk), .Q(counter[5]) );
  DFFPOSX1 counter_reg_6_ ( .D(n184), .CLK(clk), .Q(counter[6]) );
  DFFPOSX1 counter_reg_7_ ( .D(n183), .CLK(clk), .Q(counter[7]) );
  DFFPOSX1 counter_reg_8_ ( .D(n182), .CLK(clk), .Q(counter[8]) );
  DFFPOSX1 counter_reg_9_ ( .D(n181), .CLK(clk), .Q(counter[9]) );
  DFFPOSX1 counter_reg_10_ ( .D(n180), .CLK(clk), .Q(counter[10]) );
  DFFPOSX1 counter_reg_11_ ( .D(n179), .CLK(clk), .Q(counter[11]) );
  DFFPOSX1 counter_reg_12_ ( .D(n178), .CLK(clk), .Q(counter[12]) );
  DFFPOSX1 counter_reg_13_ ( .D(n177), .CLK(clk), .Q(counter[13]) );
  DFFPOSX1 counter_reg_14_ ( .D(n176), .CLK(clk), .Q(counter[14]) );
  DFFPOSX1 counter_reg_15_ ( .D(n175), .CLK(clk), .Q(counter[15]) );
  DFFPOSX1 counter_reg_16_ ( .D(n174), .CLK(clk), .Q(counter[16]) );
  DFFPOSX1 counter_reg_17_ ( .D(n173), .CLK(clk), .Q(counter[17]) );
  DFFPOSX1 counter_reg_18_ ( .D(n172), .CLK(clk), .Q(counter[18]) );
  DFFPOSX1 resetbar_reg ( .D(n30), .CLK(clk), .Q(resetbar) );
  DFFPOSX1 webar_reg ( .D(n8), .CLK(clk), .Q(webar) );
  DFFPOSX1 casbar_reg ( .D(n28), .CLK(clk), .Q(casbar) );
  DFFPOSX1 rasbar_reg ( .D(n29), .CLK(clk), .Q(rasbar) );
  DFFPOSX1 ready_reg ( .D(n171), .CLK(clk), .Q(ready) );
  DFFPOSX1 cke_reg ( .D(n31), .CLK(clk), .Q(cke) );
  DFFPOSX1 a_reg_10_ ( .D(n165), .CLK(clk), .Q(a[10]) );
  DFFPOSX1 a_reg_8_ ( .D(n32), .CLK(clk), .Q(a[8]) );
  DFFPOSX1 a_reg_4_ ( .D(n6), .CLK(clk), .Q(a[4]) );
  DFFPOSX1 ba_reg_1_ ( .D(n254), .CLK(clk), .Q(ba[1]) );
  DFFPOSX1 ba_reg_0_ ( .D(n7), .CLK(clk), .Q(ba[0]) );
  NAND3X1 U61 ( .A(n195), .B(n50), .C(n52), .Y(n162) );
  NAND3X1 U63 ( .A(counter[3]), .B(n271), .C(n234), .Y(n60) );
  AOI22X1 U64 ( .A(n65), .B(n234), .C(ba[1]), .D(n241), .Y(n64) );
  NAND3X1 U65 ( .A(n192), .B(n195), .C(n51), .Y(n163) );
  OAI21X1 U72 ( .A(n245), .B(n71), .C(n219), .Y(n165) );
  OAI21X1 U74 ( .A(n261), .B(n260), .C(n73), .Y(n71) );
  OAI21X1 U75 ( .A(n233), .B(n228), .C(n241), .Y(n73) );
  NAND3X1 U77 ( .A(n70), .B(n215), .C(n265), .Y(n78) );
  OAI21X1 U80 ( .A(n81), .B(n265), .C(n255), .Y(n80) );
  NOR3X1 U81 ( .A(n216), .B(n267), .C(n242), .Y(n81) );
  NAND3X1 U84 ( .A(n70), .B(n87), .C(n88), .Y(n86) );
  OAI21X1 U86 ( .A(n49), .B(n233), .C(n257), .Y(n87) );
  AOI21X1 U87 ( .A(n90), .B(n91), .C(n88), .Y(n89) );
  NOR3X1 U88 ( .A(n242), .B(n262), .C(n220), .Y(n88) );
  NAND3X1 U90 ( .A(n93), .B(n94), .C(n95), .Y(n84) );
  NOR3X1 U91 ( .A(n54), .B(n239), .C(n231), .Y(n95) );
  NAND3X1 U93 ( .A(n285), .B(n286), .C(n280), .Y(n96) );
  NOR3X1 U94 ( .A(n224), .B(counter[10]), .C(n281), .Y(n94) );
  NOR3X1 U96 ( .A(n284), .B(n273), .C(n282), .Y(n93) );
  NOR3X1 U97 ( .A(n213), .B(n239), .C(n225), .Y(n91) );
  NAND3X1 U100 ( .A(n284), .B(n285), .C(n214), .Y(n100) );
  NOR3X1 U102 ( .A(n53), .B(n55), .C(n56), .Y(n90) );
  NAND3X1 U105 ( .A(n278), .B(n279), .C(n106), .Y(n103) );
  NAND3X1 U110 ( .A(n221), .B(n110), .C(n70), .Y(n107) );
  NAND3X1 U112 ( .A(n48), .B(n221), .C(n70), .Y(n112) );
  NAND3X1 U113 ( .A(n114), .B(n193), .C(n263), .Y(n113) );
  NAND3X1 U114 ( .A(n194), .B(n82), .C(n199), .Y(n116) );
  OAI21X1 U116 ( .A(n227), .B(n245), .C(n226), .Y(n171) );
  AOI21X1 U118 ( .A(n255), .B(n264), .C(RESET), .Y(n119) );
  OAI21X1 U119 ( .A(n248), .B(n286), .C(n230), .Y(n172) );
  OAI21X1 U121 ( .A(n248), .B(n285), .C(n223), .Y(n173) );
  OAI21X1 U123 ( .A(n250), .B(n284), .C(n218), .Y(n174) );
  OAI21X1 U125 ( .A(n249), .B(n283), .C(n212), .Y(n175) );
  OAI21X1 U127 ( .A(n249), .B(n282), .C(n210), .Y(n176) );
  OAI21X1 U129 ( .A(n248), .B(n281), .C(n208), .Y(n177) );
  OAI21X1 U131 ( .A(n250), .B(n280), .C(n206), .Y(n178) );
  OAI21X1 U133 ( .A(n250), .B(n279), .C(n204), .Y(n179) );
  OAI21X1 U135 ( .A(n249), .B(n278), .C(n202), .Y(n180) );
  OAI21X1 U137 ( .A(n248), .B(n277), .C(n217), .Y(n181) );
  OAI21X1 U139 ( .A(n248), .B(n275), .C(n211), .Y(n182) );
  OAI21X1 U141 ( .A(n250), .B(n274), .C(n229), .Y(n183) );
  OAI21X1 U143 ( .A(n249), .B(n273), .C(n222), .Y(n184) );
  OAI21X1 U145 ( .A(n249), .B(n272), .C(n207), .Y(n185) );
  OAI21X1 U147 ( .A(n248), .B(n270), .C(n209), .Y(n186) );
  OAI21X1 U149 ( .A(n250), .B(n267), .C(n201), .Y(n187) );
  OAI21X1 U151 ( .A(n250), .B(n266), .C(n200), .Y(n188) );
  OAI21X1 U153 ( .A(n249), .B(n262), .C(n205), .Y(n189) );
  OAI21X1 U155 ( .A(n248), .B(n259), .C(n203), .Y(n190) );
  OAI21X1 U157 ( .A(RESET), .B(n240), .C(n245), .Y(n191) );
  OAI21X1 U160 ( .A(n110), .B(n196), .C(n255), .Y(n142) );
  NAND3X1 U161 ( .A(n193), .B(n194), .C(n114), .Y(n145) );
  NAND3X1 U162 ( .A(n243), .B(n268), .C(counter[12]), .Y(n147) );
  NAND3X1 U163 ( .A(n278), .B(n279), .C(n235), .Y(n146) );
  NAND3X1 U165 ( .A(n268), .B(n276), .C(n243), .Y(n115) );
  NAND3X1 U166 ( .A(n82), .B(n228), .C(n199), .Y(n144) );
  NAND3X1 U169 ( .A(n244), .B(n276), .C(n268), .Y(n75) );
  NAND3X1 U170 ( .A(n106), .B(counter[3]), .C(counter[7]), .Y(n151) );
  NAND3X1 U171 ( .A(n106), .B(counter[1]), .C(counter[2]), .Y(n153) );
  NOR3X1 U172 ( .A(counter[5]), .B(counter[6]), .C(counter[4]), .Y(n106) );
  NAND3X1 U173 ( .A(n267), .B(n274), .C(n276), .Y(n152) );
  AOI21X1 U174 ( .A(n196), .B(n255), .C(RESET), .Y(n62) );
  NAND3X1 U175 ( .A(n259), .B(n277), .C(n70), .Y(n74) );
  NAND3X1 U178 ( .A(n269), .B(n244), .C(counter[3]), .Y(n76) );
  NAND3X1 U180 ( .A(n156), .B(n272), .C(counter[4]), .Y(n155) );
  NAND3X1 U181 ( .A(n244), .B(n267), .C(n269), .Y(n68) );
  NAND3X1 U182 ( .A(n156), .B(n270), .C(counter[5]), .Y(n157) );
  NOR3X1 U183 ( .A(n232), .B(counter[7]), .C(n273), .Y(n156) );
  NAND3X1 U184 ( .A(counter[11]), .B(counter[10]), .C(n158), .Y(n154) );
  NAND3X1 U186 ( .A(counter[18]), .B(counter[17]), .C(counter[8]), .Y(n160) );
  NAND3X1 U187 ( .A(counter[15]), .B(counter[13]), .C(n238), .Y(n159) );
  ddr3_init_engine_DW01_inc_0 add_95 ( .A(counter), .SUM({n27, n26, n25, n24, 
        n23, n22, n21, n20, n19, n18, n17, n16, n15, n14, n13, n12, n11, n10, 
        n9}) );
  OR2X1 U17 ( .A(n236), .B(n237), .Y(n149) );
  OR2X1 U18 ( .A(n42), .B(n45), .Y(n82) );
  OR2X1 U19 ( .A(n43), .B(n47), .Y(n110) );
  OR2X1 U20 ( .A(n44), .B(n46), .Y(n114) );
  AND2X1 U21 ( .A(n250), .B(n240), .Y(n122) );
  AND2X1 U22 ( .A(ready), .B(n227), .Y(n120) );
  BUFX2 U23 ( .A(n64), .Y(n1) );
  BUFX2 U24 ( .A(n157), .Y(n2) );
  BUFX2 U25 ( .A(n155), .Y(n3) );
  BUFX2 U26 ( .A(n151), .Y(n4) );
  BUFX2 U27 ( .A(n116), .Y(n5) );
  OR2X1 U28 ( .A(n197), .B(n198), .Y(n196) );
  OR2X1 U29 ( .A(n260), .B(n65), .Y(n198) );
  BUFX2 U30 ( .A(n163), .Y(n6) );
  BUFX2 U31 ( .A(n162), .Y(n7) );
  AND2X1 U32 ( .A(n39), .B(n33), .Y(n170) );
  INVX1 U33 ( .A(n170), .Y(n8) );
  AND2X1 U34 ( .A(n143), .B(n36), .Y(n169) );
  INVX1 U35 ( .A(n169), .Y(n28) );
  AND2X1 U36 ( .A(n143), .B(n37), .Y(n168) );
  INVX1 U37 ( .A(n168), .Y(n29) );
  AND2X1 U38 ( .A(n40), .B(n34), .Y(n167) );
  INVX1 U39 ( .A(n167), .Y(n30) );
  AND2X1 U40 ( .A(n41), .B(n35), .Y(n166) );
  INVX1 U41 ( .A(n166), .Y(n31) );
  AND2X1 U42 ( .A(n192), .B(n38), .Y(n164) );
  INVX1 U43 ( .A(n164), .Y(n32) );
  BUFX2 U44 ( .A(n112), .Y(n33) );
  BUFX2 U45 ( .A(n86), .Y(n34) );
  BUFX2 U46 ( .A(n78), .Y(n35) );
  AND2X1 U47 ( .A(casbar), .B(n346), .Y(n109) );
  INVX1 U48 ( .A(n109), .Y(n36) );
  AND2X1 U49 ( .A(rasbar), .B(n346), .Y(n108) );
  INVX1 U50 ( .A(n108), .Y(n37) );
  AND2X1 U51 ( .A(a[8]), .B(n241), .Y(n69) );
  INVX1 U52 ( .A(n69), .Y(n38) );
  AND2X1 U53 ( .A(webar), .B(n346), .Y(n111) );
  INVX1 U54 ( .A(n111), .Y(n39) );
  AND2X1 U55 ( .A(resetbar), .B(n256), .Y(n85) );
  INVX1 U56 ( .A(n85), .Y(n40) );
  AND2X1 U57 ( .A(cke), .B(n79), .Y(n77) );
  INVX1 U58 ( .A(n77), .Y(n41) );
  BUFX2 U59 ( .A(n152), .Y(n42) );
  BUFX2 U60 ( .A(n144), .Y(n43) );
  BUFX2 U62 ( .A(n146), .Y(n44) );
  BUFX2 U66 ( .A(n153), .Y(n45) );
  BUFX2 U67 ( .A(n147), .Y(n46) );
  BUFX2 U68 ( .A(n145), .Y(n47) );
  BUFX2 U69 ( .A(n113), .Y(n48) );
  BUFX2 U70 ( .A(n89), .Y(n49) );
  BUFX2 U71 ( .A(n60), .Y(n50) );
  AND2X1 U73 ( .A(a[4]), .B(n241), .Y(n67) );
  INVX1 U76 ( .A(n67), .Y(n51) );
  AND2X1 U78 ( .A(ba[0]), .B(n241), .Y(n61) );
  INVX1 U79 ( .A(n61), .Y(n52) );
  BUFX2 U82 ( .A(n103), .Y(n53) );
  BUFX2 U83 ( .A(n96), .Y(n54) );
  AND2X1 U85 ( .A(n282), .B(n283), .Y(n104) );
  INVX1 U89 ( .A(n104), .Y(n55) );
  AND2X1 U92 ( .A(n280), .B(n281), .Y(n105) );
  INVX1 U95 ( .A(n105), .Y(n56) );
  BUFX2 U98 ( .A(n68), .Y(n57) );
  BUFX2 U99 ( .A(n76), .Y(n58) );
  AND2X1 U101 ( .A(n271), .B(n244), .Y(n65) );
  BUFX2 U103 ( .A(n107), .Y(n143) );
  AND2X1 U104 ( .A(n260), .B(n234), .Y(n66) );
  INVX1 U106 ( .A(n66), .Y(n192) );
  BUFX2 U107 ( .A(n115), .Y(n193) );
  AND2X1 U108 ( .A(n243), .B(n269), .Y(n117) );
  INVX1 U109 ( .A(n117), .Y(n194) );
  AND2X1 U111 ( .A(n197), .B(n234), .Y(n59) );
  INVX1 U115 ( .A(n59), .Y(n195) );
  INVX1 U117 ( .A(n57), .Y(n197) );
  AND2X1 U120 ( .A(n243), .B(n271), .Y(n118) );
  INVX1 U122 ( .A(n118), .Y(n199) );
  AND2X1 U124 ( .A(n11), .B(n251), .Y(n138) );
  INVX1 U126 ( .A(n138), .Y(n200) );
  AND2X1 U128 ( .A(n12), .B(n251), .Y(n137) );
  INVX1 U130 ( .A(n137), .Y(n201) );
  AND2X1 U132 ( .A(n19), .B(n252), .Y(n130) );
  INVX1 U134 ( .A(n130), .Y(n202) );
  AND2X1 U136 ( .A(n9), .B(n251), .Y(n140) );
  INVX1 U138 ( .A(n140), .Y(n203) );
  AND2X1 U140 ( .A(n20), .B(n252), .Y(n129) );
  INVX1 U142 ( .A(n129), .Y(n204) );
  AND2X1 U144 ( .A(n10), .B(n251), .Y(n139) );
  INVX1 U146 ( .A(n139), .Y(n205) );
  AND2X1 U148 ( .A(n21), .B(n252), .Y(n128) );
  INVX1 U150 ( .A(n128), .Y(n206) );
  AND2X1 U152 ( .A(n14), .B(n251), .Y(n135) );
  INVX1 U154 ( .A(n135), .Y(n207) );
  AND2X1 U156 ( .A(n22), .B(n252), .Y(n127) );
  INVX1 U158 ( .A(n127), .Y(n208) );
  AND2X1 U159 ( .A(n13), .B(n251), .Y(n136) );
  INVX1 U164 ( .A(n136), .Y(n209) );
  AND2X1 U167 ( .A(n23), .B(n252), .Y(n126) );
  INVX1 U168 ( .A(n126), .Y(n210) );
  AND2X1 U176 ( .A(n17), .B(n251), .Y(n132) );
  INVX1 U177 ( .A(n132), .Y(n211) );
  AND2X1 U179 ( .A(n24), .B(n252), .Y(n125) );
  INVX1 U185 ( .A(n125), .Y(n212) );
  BUFX2 U188 ( .A(n100), .Y(n213) );
  OR2X1 U189 ( .A(counter[1]), .B(counter[18]), .Y(n102) );
  INVX1 U190 ( .A(n102), .Y(n214) );
  AND2X1 U191 ( .A(n257), .B(n80), .Y(n79) );
  INVX1 U192 ( .A(n79), .Y(n215) );
  AND2X1 U193 ( .A(n262), .B(n270), .Y(n83) );
  INVX1 U194 ( .A(n83), .Y(n216) );
  AND2X1 U195 ( .A(n18), .B(n251), .Y(n131) );
  INVX1 U196 ( .A(n131), .Y(n217) );
  AND2X1 U197 ( .A(n25), .B(n252), .Y(n124) );
  INVX1 U198 ( .A(n124), .Y(n218) );
  AND2X1 U199 ( .A(a[10]), .B(n253), .Y(n72) );
  INVX1 U200 ( .A(n72), .Y(n219) );
  AND2X1 U201 ( .A(n267), .B(counter[4]), .Y(n92) );
  INVX1 U202 ( .A(n92), .Y(n220) );
  AND2X1 U203 ( .A(n257), .B(n142), .Y(n346) );
  INVX1 U204 ( .A(n346), .Y(n221) );
  AND2X1 U205 ( .A(n15), .B(n251), .Y(n134) );
  INVX1 U206 ( .A(n134), .Y(n222) );
  AND2X1 U207 ( .A(n26), .B(n252), .Y(n123) );
  INVX1 U208 ( .A(n123), .Y(n223) );
  AND2X1 U209 ( .A(counter[11]), .B(counter[15]), .Y(n99) );
  INVX1 U210 ( .A(n99), .Y(n224) );
  AND2X1 U211 ( .A(n266), .B(n267), .Y(n101) );
  INVX1 U212 ( .A(n101), .Y(n225) );
  INVX1 U213 ( .A(n120), .Y(n226) );
  BUFX2 U214 ( .A(n119), .Y(n227) );
  BUFX2 U215 ( .A(n75), .Y(n228) );
  AND2X1 U216 ( .A(n16), .B(n251), .Y(n133) );
  INVX1 U217 ( .A(n133), .Y(n229) );
  AND2X1 U218 ( .A(n27), .B(n252), .Y(n121) );
  INVX1 U219 ( .A(n121), .Y(n230) );
  AND2X1 U220 ( .A(n266), .B(n272), .Y(n98) );
  INVX1 U221 ( .A(n98), .Y(n231) );
  BUFX2 U222 ( .A(n154), .Y(n232) );
  AND2X1 U223 ( .A(n280), .B(n235), .Y(n158) );
  BUFX2 U224 ( .A(n74), .Y(n233) );
  OR2X1 U225 ( .A(n245), .B(n241), .Y(n63) );
  INVX1 U226 ( .A(n63), .Y(n234) );
  INVX1 U227 ( .A(n149), .Y(n235) );
  BUFX2 U228 ( .A(n159), .Y(n236) );
  BUFX2 U229 ( .A(n160), .Y(n237) );
  OR2X1 U230 ( .A(counter[16]), .B(counter[14]), .Y(n161) );
  INVX1 U231 ( .A(n161), .Y(n238) );
  AND2X1 U232 ( .A(n274), .B(n275), .Y(n97) );
  INVX1 U233 ( .A(n97), .Y(n239) );
  AND2X1 U234 ( .A(INIT), .B(n258), .Y(n141) );
  INVX1 U235 ( .A(n141), .Y(n240) );
  BUFX2 U236 ( .A(n62), .Y(n241) );
  BUFX2 U237 ( .A(n84), .Y(n242) );
  OR2X1 U238 ( .A(n266), .B(counter[1]), .Y(n148) );
  INVX1 U239 ( .A(n148), .Y(n243) );
  OR2X1 U240 ( .A(n262), .B(counter[2]), .Y(n150) );
  INVX1 U241 ( .A(n150), .Y(n244) );
  AND2X1 U242 ( .A(flag), .B(n257), .Y(n70) );
  INVX1 U243 ( .A(n70), .Y(n245) );
  INVX1 U244 ( .A(n233), .Y(n255) );
  BUFX2 U245 ( .A(n122), .Y(n251) );
  BUFX2 U246 ( .A(n122), .Y(n252) );
  INVX1 U247 ( .A(n228), .Y(n261) );
  INVX1 U248 ( .A(n232), .Y(n276) );
  INVX1 U249 ( .A(n58), .Y(n260) );
  INVX1 U250 ( .A(n5), .Y(n263) );
  INVX1 U251 ( .A(n82), .Y(n265) );
  INVX1 U252 ( .A(n1), .Y(n254) );
  INVX1 U253 ( .A(n3), .Y(n271) );
  INVX1 U254 ( .A(n2), .Y(n269) );
  INVX1 U255 ( .A(n73), .Y(n253) );
  INVX1 U256 ( .A(counter[12]), .Y(n280) );
  INVX1 U257 ( .A(flag), .Y(n258) );
  INVX1 U258 ( .A(n114), .Y(n264) );
  INVX1 U259 ( .A(counter[3]), .Y(n267) );
  INVX1 U260 ( .A(n87), .Y(n256) );
  BUFX2 U261 ( .A(n246), .Y(n248) );
  BUFX2 U262 ( .A(n247), .Y(n249) );
  BUFX2 U263 ( .A(n191), .Y(n250) );
  INVX1 U264 ( .A(counter[1]), .Y(n262) );
  INVX1 U265 ( .A(counter[2]), .Y(n266) );
  INVX1 U266 ( .A(RESET), .Y(n257) );
  INVX1 U267 ( .A(counter[4]), .Y(n270) );
  INVX1 U268 ( .A(counter[6]), .Y(n273) );
  INVX1 U269 ( .A(n4), .Y(n268) );
  INVX1 U270 ( .A(counter[11]), .Y(n279) );
  INVX1 U271 ( .A(counter[10]), .Y(n278) );
  INVX1 U272 ( .A(counter[7]), .Y(n274) );
  INVX1 U273 ( .A(counter[5]), .Y(n272) );
  INVX1 U274 ( .A(counter[16]), .Y(n284) );
  INVX1 U275 ( .A(counter[17]), .Y(n285) );
  INVX1 U276 ( .A(counter[13]), .Y(n281) );
  INVX1 U277 ( .A(counter[14]), .Y(n282) );
  INVX1 U278 ( .A(counter[18]), .Y(n286) );
  INVX1 U279 ( .A(counter[15]), .Y(n283) );
  INVX1 U280 ( .A(counter[8]), .Y(n275) );
  INVX1 U281 ( .A(counter[0]), .Y(n259) );
  INVX1 U282 ( .A(counter[9]), .Y(n277) );
  OAI21X1 U283 ( .A(RESET), .B(n240), .C(n245), .Y(n246) );
  OAI21X1 U284 ( .A(RESET), .B(n240), .C(n245), .Y(n247) );
endmodule


module ddr3_ring_buffer8 ( dout, listen, strobe, readPtr, din, reset );
  output [15:0] dout;
  input [1:0] strobe;
  input [2:0] readPtr;
  input [15:0] din;
  input listen, reset;
  wire   dStrobe0, n_0_net_, F0, dStrobe1, dStrobe2, dnStrobe, dStrobe3,
         n_1_net_, dStrobe4, dStrobe5, dpStrobe, n72, n73, n74, n76, n78, n80,
         n82, n84, n86, n88, n90, n92, n94, n96, n98, n100, n102, n104, n106,
         n108, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n315, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n448, n452, n453, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n75, n77, n79, n81, n83, n85, n87, n89, n91, n93,
         n95, n97, n99, n101, n103, n105, n107, n109, n229, n230, n231, n232,
         n314, n316, n447, n450, n451, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n465, n466, n467, n468, n469, n470, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n487, n488, n489, n490, n491, n492, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n509, n510, n511, n512, n513, n514, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n531, n532,
         n533, n534, n535, n536, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n553, n554, n555, n556,
         n557, n558, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n576, n577, n578, n579, n580,
         n581, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n601, n602, n603, n604,
         n605, n606, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n624, n625, n626, n627, n628,
         n629, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674;
  wire   [3:0] nStrobe;
  wire   [3:0] pStrobe;
  wire   [1:0] count;
  wire   [15:0] r0;
  wire   [15:0] r2;
  wire   [15:0] r4;
  wire   [15:0] r6;
  wire   [15:0] r1;
  wire   [15:0] r3;
  wire   [15:0] r5;
  wire   [15:0] r7;

  CLKBUF2 DELAY0 ( .A(n_0_net_), .Y(dStrobe0) );
  CLKBUF2 DELAY1 ( .A(dStrobe0), .Y(dStrobe1) );
  CLKBUF2 DELAY2 ( .A(dStrobe1), .Y(dStrobe2) );
  CLKBUF2 DELAY3 ( .A(dStrobe2), .Y(dnStrobe) );
  CLKBUF2 DELAYN0 ( .A(dnStrobe), .Y(nStrobe[0]) );
  CLKBUF2 DELAYN1 ( .A(dnStrobe), .Y(nStrobe[1]) );
  CLKBUF2 DELAYN2 ( .A(dnStrobe), .Y(nStrobe[2]) );
  CLKBUF2 DELAYN3 ( .A(dnStrobe), .Y(nStrobe[3]) );
  CLKBUF2 DELAY4 ( .A(n_1_net_), .Y(dStrobe3) );
  CLKBUF2 DELAY5 ( .A(dStrobe3), .Y(dStrobe4) );
  CLKBUF2 DELAY6 ( .A(dStrobe4), .Y(dStrobe5) );
  CLKBUF2 DELAY7 ( .A(dStrobe5), .Y(dpStrobe) );
  CLKBUF2 DELAYP0 ( .A(dpStrobe), .Y(pStrobe[0]) );
  CLKBUF2 DELAYP1 ( .A(dpStrobe), .Y(pStrobe[1]) );
  CLKBUF2 DELAYP2 ( .A(dpStrobe), .Y(pStrobe[2]) );
  CLKBUF2 DELAYP3 ( .A(dpStrobe), .Y(pStrobe[3]) );
  DFFSR count_reg_0_ ( .D(n453), .CLK(n651), .R(n649), .S(1'b1), .Q(count[0])
         );
  DFFSR F0_reg ( .D(n448), .CLK(n651), .R(n649), .S(n668), .Q(F0) );
  DFFSR count_reg_1_ ( .D(n452), .CLK(n651), .R(n649), .S(1'b1), .Q(count[1])
         );
  DFFPOSX1 r0_reg_15_ ( .D(n445), .CLK(pStrobe[0]), .Q(r0[15]) );
  DFFPOSX1 r0_reg_14_ ( .D(n444), .CLK(pStrobe[0]), .Q(r0[14]) );
  DFFPOSX1 r0_reg_13_ ( .D(n443), .CLK(pStrobe[0]), .Q(r0[13]) );
  DFFPOSX1 r0_reg_12_ ( .D(n442), .CLK(pStrobe[0]), .Q(r0[12]) );
  DFFPOSX1 r0_reg_11_ ( .D(n441), .CLK(pStrobe[0]), .Q(r0[11]) );
  DFFPOSX1 r0_reg_10_ ( .D(n440), .CLK(pStrobe[0]), .Q(r0[10]) );
  DFFPOSX1 r0_reg_9_ ( .D(n439), .CLK(pStrobe[0]), .Q(r0[9]) );
  DFFPOSX1 r0_reg_8_ ( .D(n438), .CLK(pStrobe[0]), .Q(r0[8]) );
  DFFPOSX1 r0_reg_7_ ( .D(n437), .CLK(pStrobe[0]), .Q(r0[7]) );
  DFFPOSX1 r0_reg_6_ ( .D(n436), .CLK(pStrobe[0]), .Q(r0[6]) );
  DFFPOSX1 r0_reg_5_ ( .D(n435), .CLK(pStrobe[0]), .Q(r0[5]) );
  DFFPOSX1 r0_reg_4_ ( .D(n434), .CLK(pStrobe[0]), .Q(r0[4]) );
  DFFPOSX1 r0_reg_3_ ( .D(n433), .CLK(pStrobe[0]), .Q(r0[3]) );
  DFFPOSX1 r0_reg_2_ ( .D(n432), .CLK(pStrobe[0]), .Q(r0[2]) );
  DFFPOSX1 r0_reg_1_ ( .D(n431), .CLK(pStrobe[0]), .Q(r0[1]) );
  DFFPOSX1 r0_reg_0_ ( .D(n430), .CLK(pStrobe[0]), .Q(r0[0]) );
  DFFPOSX1 r2_reg_15_ ( .D(n429), .CLK(pStrobe[1]), .Q(r2[15]) );
  DFFPOSX1 r2_reg_14_ ( .D(n428), .CLK(pStrobe[1]), .Q(r2[14]) );
  DFFPOSX1 r2_reg_13_ ( .D(n427), .CLK(pStrobe[1]), .Q(r2[13]) );
  DFFPOSX1 r2_reg_12_ ( .D(n426), .CLK(pStrobe[1]), .Q(r2[12]) );
  DFFPOSX1 r2_reg_11_ ( .D(n425), .CLK(pStrobe[1]), .Q(r2[11]) );
  DFFPOSX1 r2_reg_10_ ( .D(n424), .CLK(pStrobe[1]), .Q(r2[10]) );
  DFFPOSX1 r2_reg_9_ ( .D(n423), .CLK(pStrobe[1]), .Q(r2[9]) );
  DFFPOSX1 r2_reg_8_ ( .D(n422), .CLK(pStrobe[1]), .Q(r2[8]) );
  DFFPOSX1 r2_reg_7_ ( .D(n421), .CLK(pStrobe[1]), .Q(r2[7]) );
  DFFPOSX1 r2_reg_6_ ( .D(n420), .CLK(pStrobe[1]), .Q(r2[6]) );
  DFFPOSX1 r2_reg_5_ ( .D(n419), .CLK(pStrobe[1]), .Q(r2[5]) );
  DFFPOSX1 r2_reg_4_ ( .D(n418), .CLK(pStrobe[1]), .Q(r2[4]) );
  DFFPOSX1 r2_reg_3_ ( .D(n417), .CLK(pStrobe[1]), .Q(r2[3]) );
  DFFPOSX1 r2_reg_2_ ( .D(n416), .CLK(pStrobe[1]), .Q(r2[2]) );
  DFFPOSX1 r2_reg_1_ ( .D(n415), .CLK(pStrobe[1]), .Q(r2[1]) );
  DFFPOSX1 r2_reg_0_ ( .D(n414), .CLK(pStrobe[1]), .Q(r2[0]) );
  DFFPOSX1 r4_reg_15_ ( .D(n413), .CLK(pStrobe[2]), .Q(r4[15]) );
  DFFPOSX1 r4_reg_14_ ( .D(n412), .CLK(pStrobe[2]), .Q(r4[14]) );
  DFFPOSX1 r4_reg_13_ ( .D(n411), .CLK(pStrobe[2]), .Q(r4[13]) );
  DFFPOSX1 r4_reg_12_ ( .D(n410), .CLK(pStrobe[2]), .Q(r4[12]) );
  DFFPOSX1 r4_reg_11_ ( .D(n409), .CLK(pStrobe[2]), .Q(r4[11]) );
  DFFPOSX1 r4_reg_10_ ( .D(n408), .CLK(pStrobe[2]), .Q(r4[10]) );
  DFFPOSX1 r4_reg_9_ ( .D(n407), .CLK(pStrobe[2]), .Q(r4[9]) );
  DFFPOSX1 r4_reg_8_ ( .D(n406), .CLK(pStrobe[2]), .Q(r4[8]) );
  DFFPOSX1 r4_reg_7_ ( .D(n405), .CLK(pStrobe[2]), .Q(r4[7]) );
  DFFPOSX1 r4_reg_6_ ( .D(n404), .CLK(pStrobe[2]), .Q(r4[6]) );
  DFFPOSX1 r4_reg_5_ ( .D(n403), .CLK(pStrobe[2]), .Q(r4[5]) );
  DFFPOSX1 r4_reg_4_ ( .D(n402), .CLK(pStrobe[2]), .Q(r4[4]) );
  DFFPOSX1 r4_reg_3_ ( .D(n401), .CLK(pStrobe[2]), .Q(r4[3]) );
  DFFPOSX1 r4_reg_2_ ( .D(n400), .CLK(pStrobe[2]), .Q(r4[2]) );
  DFFPOSX1 r4_reg_1_ ( .D(n399), .CLK(pStrobe[2]), .Q(r4[1]) );
  DFFPOSX1 r4_reg_0_ ( .D(n398), .CLK(pStrobe[2]), .Q(r4[0]) );
  DFFPOSX1 r6_reg_15_ ( .D(n397), .CLK(pStrobe[3]), .Q(r6[15]) );
  DFFPOSX1 r6_reg_14_ ( .D(n396), .CLK(pStrobe[3]), .Q(r6[14]) );
  DFFPOSX1 r6_reg_13_ ( .D(n395), .CLK(pStrobe[3]), .Q(r6[13]) );
  DFFPOSX1 r6_reg_12_ ( .D(n394), .CLK(pStrobe[3]), .Q(r6[12]) );
  DFFPOSX1 r6_reg_11_ ( .D(n393), .CLK(pStrobe[3]), .Q(r6[11]) );
  DFFPOSX1 r6_reg_10_ ( .D(n392), .CLK(pStrobe[3]), .Q(r6[10]) );
  DFFPOSX1 r6_reg_9_ ( .D(n391), .CLK(pStrobe[3]), .Q(r6[9]) );
  DFFPOSX1 r6_reg_8_ ( .D(n390), .CLK(pStrobe[3]), .Q(r6[8]) );
  DFFPOSX1 r6_reg_7_ ( .D(n389), .CLK(pStrobe[3]), .Q(r6[7]) );
  DFFPOSX1 r6_reg_6_ ( .D(n388), .CLK(pStrobe[3]), .Q(r6[6]) );
  DFFPOSX1 r6_reg_5_ ( .D(n387), .CLK(pStrobe[3]), .Q(r6[5]) );
  DFFPOSX1 r6_reg_4_ ( .D(n386), .CLK(pStrobe[3]), .Q(r6[4]) );
  DFFPOSX1 r6_reg_3_ ( .D(n385), .CLK(pStrobe[3]), .Q(r6[3]) );
  DFFPOSX1 r6_reg_2_ ( .D(n384), .CLK(pStrobe[3]), .Q(r6[2]) );
  DFFPOSX1 r6_reg_1_ ( .D(n383), .CLK(pStrobe[3]), .Q(r6[1]) );
  DFFPOSX1 r6_reg_0_ ( .D(n382), .CLK(pStrobe[3]), .Q(r6[0]) );
  DFFNEGX1 r1_reg_15_ ( .D(n381), .CLK(nStrobe[0]), .Q(r1[15]) );
  DFFNEGX1 r1_reg_14_ ( .D(n380), .CLK(nStrobe[0]), .Q(r1[14]) );
  DFFNEGX1 r1_reg_13_ ( .D(n379), .CLK(nStrobe[0]), .Q(r1[13]) );
  DFFNEGX1 r1_reg_12_ ( .D(n378), .CLK(nStrobe[0]), .Q(r1[12]) );
  DFFNEGX1 r1_reg_11_ ( .D(n377), .CLK(nStrobe[0]), .Q(r1[11]) );
  DFFNEGX1 r1_reg_10_ ( .D(n376), .CLK(nStrobe[0]), .Q(r1[10]) );
  DFFNEGX1 r1_reg_9_ ( .D(n375), .CLK(nStrobe[0]), .Q(r1[9]) );
  DFFNEGX1 r1_reg_8_ ( .D(n374), .CLK(nStrobe[0]), .Q(r1[8]) );
  DFFNEGX1 r1_reg_7_ ( .D(n373), .CLK(nStrobe[0]), .Q(r1[7]) );
  DFFNEGX1 r1_reg_6_ ( .D(n372), .CLK(nStrobe[0]), .Q(r1[6]) );
  DFFNEGX1 r1_reg_5_ ( .D(n371), .CLK(nStrobe[0]), .Q(r1[5]) );
  DFFNEGX1 r1_reg_4_ ( .D(n370), .CLK(nStrobe[0]), .Q(r1[4]) );
  DFFNEGX1 r1_reg_3_ ( .D(n369), .CLK(nStrobe[0]), .Q(r1[3]) );
  DFFNEGX1 r1_reg_2_ ( .D(n368), .CLK(nStrobe[0]), .Q(r1[2]) );
  DFFNEGX1 r1_reg_1_ ( .D(n367), .CLK(nStrobe[0]), .Q(r1[1]) );
  DFFNEGX1 r1_reg_0_ ( .D(n366), .CLK(nStrobe[0]), .Q(r1[0]) );
  DFFNEGX1 r3_reg_15_ ( .D(n365), .CLK(nStrobe[1]), .Q(r3[15]) );
  DFFNEGX1 r3_reg_14_ ( .D(n364), .CLK(nStrobe[1]), .Q(r3[14]) );
  DFFNEGX1 r3_reg_13_ ( .D(n363), .CLK(nStrobe[1]), .Q(r3[13]) );
  DFFNEGX1 r3_reg_12_ ( .D(n362), .CLK(nStrobe[1]), .Q(r3[12]) );
  DFFNEGX1 r3_reg_11_ ( .D(n361), .CLK(nStrobe[1]), .Q(r3[11]) );
  DFFNEGX1 r3_reg_10_ ( .D(n360), .CLK(nStrobe[1]), .Q(r3[10]) );
  DFFNEGX1 r3_reg_9_ ( .D(n359), .CLK(nStrobe[1]), .Q(r3[9]) );
  DFFNEGX1 r3_reg_8_ ( .D(n358), .CLK(nStrobe[1]), .Q(r3[8]) );
  DFFNEGX1 r3_reg_7_ ( .D(n357), .CLK(nStrobe[1]), .Q(r3[7]) );
  DFFNEGX1 r3_reg_6_ ( .D(n356), .CLK(nStrobe[1]), .Q(r3[6]) );
  DFFNEGX1 r3_reg_5_ ( .D(n355), .CLK(nStrobe[1]), .Q(r3[5]) );
  DFFNEGX1 r3_reg_4_ ( .D(n354), .CLK(nStrobe[1]), .Q(r3[4]) );
  DFFNEGX1 r3_reg_3_ ( .D(n353), .CLK(nStrobe[1]), .Q(r3[3]) );
  DFFNEGX1 r3_reg_2_ ( .D(n352), .CLK(nStrobe[1]), .Q(r3[2]) );
  DFFNEGX1 r3_reg_1_ ( .D(n351), .CLK(nStrobe[1]), .Q(r3[1]) );
  DFFNEGX1 r3_reg_0_ ( .D(n350), .CLK(nStrobe[1]), .Q(r3[0]) );
  DFFNEGX1 r5_reg_15_ ( .D(n349), .CLK(nStrobe[2]), .Q(r5[15]) );
  DFFNEGX1 r5_reg_14_ ( .D(n348), .CLK(nStrobe[2]), .Q(r5[14]) );
  DFFNEGX1 r5_reg_13_ ( .D(n347), .CLK(nStrobe[2]), .Q(r5[13]) );
  DFFNEGX1 r5_reg_12_ ( .D(n346), .CLK(nStrobe[2]), .Q(r5[12]) );
  DFFNEGX1 r5_reg_11_ ( .D(n345), .CLK(nStrobe[2]), .Q(r5[11]) );
  DFFNEGX1 r5_reg_10_ ( .D(n344), .CLK(nStrobe[2]), .Q(r5[10]) );
  DFFNEGX1 r5_reg_9_ ( .D(n343), .CLK(nStrobe[2]), .Q(r5[9]) );
  DFFNEGX1 r5_reg_8_ ( .D(n342), .CLK(nStrobe[2]), .Q(r5[8]) );
  DFFNEGX1 r5_reg_7_ ( .D(n341), .CLK(nStrobe[2]), .Q(r5[7]) );
  DFFNEGX1 r5_reg_6_ ( .D(n340), .CLK(nStrobe[2]), .Q(r5[6]) );
  DFFNEGX1 r5_reg_5_ ( .D(n339), .CLK(nStrobe[2]), .Q(r5[5]) );
  DFFNEGX1 r5_reg_4_ ( .D(n338), .CLK(nStrobe[2]), .Q(r5[4]) );
  DFFNEGX1 r5_reg_3_ ( .D(n337), .CLK(nStrobe[2]), .Q(r5[3]) );
  DFFNEGX1 r5_reg_2_ ( .D(n336), .CLK(nStrobe[2]), .Q(r5[2]) );
  DFFNEGX1 r5_reg_1_ ( .D(n335), .CLK(nStrobe[2]), .Q(r5[1]) );
  DFFNEGX1 r5_reg_0_ ( .D(n334), .CLK(nStrobe[2]), .Q(r5[0]) );
  DFFNEGX1 r7_reg_15_ ( .D(n333), .CLK(nStrobe[3]), .Q(r7[15]) );
  DFFNEGX1 r7_reg_14_ ( .D(n332), .CLK(nStrobe[3]), .Q(r7[14]) );
  DFFNEGX1 r7_reg_13_ ( .D(n331), .CLK(nStrobe[3]), .Q(r7[13]) );
  DFFNEGX1 r7_reg_12_ ( .D(n330), .CLK(nStrobe[3]), .Q(r7[12]) );
  DFFNEGX1 r7_reg_11_ ( .D(n329), .CLK(nStrobe[3]), .Q(r7[11]) );
  DFFNEGX1 r7_reg_10_ ( .D(n328), .CLK(nStrobe[3]), .Q(r7[10]) );
  DFFNEGX1 r7_reg_9_ ( .D(n327), .CLK(nStrobe[3]), .Q(r7[9]) );
  DFFNEGX1 r7_reg_8_ ( .D(n326), .CLK(nStrobe[3]), .Q(r7[8]) );
  DFFNEGX1 r7_reg_7_ ( .D(n325), .CLK(nStrobe[3]), .Q(r7[7]) );
  DFFNEGX1 r7_reg_6_ ( .D(n324), .CLK(nStrobe[3]), .Q(r7[6]) );
  DFFNEGX1 r7_reg_5_ ( .D(n323), .CLK(nStrobe[3]), .Q(r7[5]) );
  DFFNEGX1 r7_reg_4_ ( .D(n322), .CLK(nStrobe[3]), .Q(r7[4]) );
  DFFNEGX1 r7_reg_3_ ( .D(n321), .CLK(nStrobe[3]), .Q(r7[3]) );
  DFFNEGX1 r7_reg_2_ ( .D(n320), .CLK(nStrobe[3]), .Q(r7[2]) );
  DFFNEGX1 r7_reg_1_ ( .D(n319), .CLK(nStrobe[3]), .Q(r7[1]) );
  DFFNEGX1 r7_reg_0_ ( .D(n318), .CLK(nStrobe[3]), .Q(r7[0]) );
  OAI21X1 U3 ( .A(n72), .B(n647), .C(n38), .Y(n452) );
  AOI21X1 U4 ( .A(n72), .B(n622), .C(n76), .Y(n74) );
  XOR2X1 U6 ( .A(n72), .B(n650), .Y(n453) );
  OAI21X1 U8 ( .A(n645), .B(n652), .C(n621), .Y(n318) );
  OAI21X1 U10 ( .A(n645), .B(n653), .C(n598), .Y(n319) );
  OAI21X1 U12 ( .A(n645), .B(n654), .C(n573), .Y(n320) );
  OAI21X1 U14 ( .A(n645), .B(n655), .C(n551), .Y(n321) );
  OAI21X1 U16 ( .A(n645), .B(n656), .C(n529), .Y(n322) );
  OAI21X1 U18 ( .A(n645), .B(n657), .C(n620), .Y(n323) );
  OAI21X1 U20 ( .A(n645), .B(n658), .C(n507), .Y(n324) );
  OAI21X1 U22 ( .A(n645), .B(n659), .C(n485), .Y(n325) );
  OAI21X1 U24 ( .A(n645), .B(n660), .C(n463), .Y(n326) );
  OAI21X1 U26 ( .A(n645), .B(n661), .C(n456), .Y(n327) );
  OAI21X1 U28 ( .A(n645), .B(n662), .C(n597), .Y(n328) );
  OAI21X1 U30 ( .A(n645), .B(n663), .C(n231), .Y(n329) );
  OAI21X1 U32 ( .A(n645), .B(n664), .C(n99), .Y(n330) );
  OAI21X1 U34 ( .A(n645), .B(n665), .C(n85), .Y(n331) );
  OAI21X1 U36 ( .A(n645), .B(n666), .C(n572), .Y(n332) );
  OAI21X1 U38 ( .A(n645), .B(n667), .C(n71), .Y(n333) );
  OAI21X1 U40 ( .A(n652), .B(n646), .C(n596), .Y(n334) );
  OAI21X1 U42 ( .A(n653), .B(n646), .C(n619), .Y(n335) );
  OAI21X1 U44 ( .A(n654), .B(n646), .C(n550), .Y(n336) );
  OAI21X1 U46 ( .A(n655), .B(n646), .C(n571), .Y(n337) );
  OAI21X1 U48 ( .A(n656), .B(n646), .C(n506), .Y(n338) );
  OAI21X1 U50 ( .A(n657), .B(n646), .C(n528), .Y(n339) );
  OAI21X1 U52 ( .A(n658), .B(n646), .C(n595), .Y(n340) );
  OAI21X1 U54 ( .A(n659), .B(n646), .C(n462), .Y(n341) );
  OAI21X1 U56 ( .A(n660), .B(n646), .C(n484), .Y(n342) );
  OAI21X1 U58 ( .A(n661), .B(n646), .C(n230), .Y(n343) );
  OAI21X1 U60 ( .A(n662), .B(n646), .C(n455), .Y(n344) );
  OAI21X1 U62 ( .A(n663), .B(n646), .C(n97), .Y(n345) );
  OAI21X1 U64 ( .A(n664), .B(n646), .C(n83), .Y(n346) );
  OAI21X1 U66 ( .A(n665), .B(n646), .C(n618), .Y(n347) );
  OAI21X1 U68 ( .A(n666), .B(n646), .C(n549), .Y(n348) );
  OAI21X1 U70 ( .A(n667), .B(n646), .C(n570), .Y(n349) );
  OAI21X1 U72 ( .A(n647), .B(n652), .C(n569), .Y(n350) );
  OAI21X1 U74 ( .A(n647), .B(n653), .C(n548), .Y(n351) );
  OAI21X1 U76 ( .A(n73), .B(n654), .C(n617), .Y(n352) );
  OAI21X1 U78 ( .A(n73), .B(n655), .C(n594), .Y(n353) );
  OAI21X1 U80 ( .A(n73), .B(n656), .C(n483), .Y(n354) );
  OAI21X1 U82 ( .A(n73), .B(n657), .C(n505), .Y(n355) );
  OAI21X1 U84 ( .A(n73), .B(n658), .C(n527), .Y(n356) );
  OAI21X1 U86 ( .A(n73), .B(n659), .C(n616), .Y(n357) );
  OAI21X1 U88 ( .A(n73), .B(n660), .C(n454), .Y(n358) );
  OAI21X1 U90 ( .A(n73), .B(n661), .C(n568), .Y(n359) );
  OAI21X1 U92 ( .A(n73), .B(n662), .C(n526), .Y(n360) );
  OAI21X1 U94 ( .A(n73), .B(n663), .C(n593), .Y(n361) );
  OAI21X1 U96 ( .A(n73), .B(n664), .C(n547), .Y(n362) );
  OAI21X1 U98 ( .A(n73), .B(n665), .C(n504), .Y(n363) );
  OAI21X1 U100 ( .A(n73), .B(n666), .C(n482), .Y(n364) );
  OAI21X1 U102 ( .A(n647), .B(n667), .C(n461), .Y(n365) );
  OAI21X1 U104 ( .A(n652), .B(n5), .C(n546), .Y(n366) );
  OAI21X1 U106 ( .A(n653), .B(n5), .C(n567), .Y(n367) );
  OAI21X1 U108 ( .A(n654), .B(n5), .C(n592), .Y(n368) );
  OAI21X1 U110 ( .A(n655), .B(n5), .C(n615), .Y(n369) );
  OAI21X1 U112 ( .A(n656), .B(n5), .C(n460), .Y(n370) );
  OAI21X1 U114 ( .A(n657), .B(n5), .C(n545), .Y(n371) );
  OAI21X1 U116 ( .A(n658), .B(n5), .C(n451), .Y(n372) );
  OAI21X1 U118 ( .A(n659), .B(n5), .C(n525), .Y(n373) );
  OAI21X1 U120 ( .A(n660), .B(n5), .C(n503), .Y(n374) );
  OAI21X1 U122 ( .A(n661), .B(n5), .C(n481), .Y(n375) );
  OAI21X1 U124 ( .A(n662), .B(n5), .C(n229), .Y(n376) );
  OAI21X1 U126 ( .A(n663), .B(n5), .C(n81), .Y(n377) );
  OAI21X1 U128 ( .A(n664), .B(n5), .C(n70), .Y(n378) );
  OAI21X1 U130 ( .A(n665), .B(n5), .C(n591), .Y(n379) );
  OAI21X1 U132 ( .A(n666), .B(n5), .C(n614), .Y(n380) );
  OAI21X1 U134 ( .A(n667), .B(n5), .C(n524), .Y(n381) );
  OAI21X1 U136 ( .A(n645), .B(n652), .C(n65), .Y(n382) );
  OAI21X1 U138 ( .A(n645), .B(n653), .C(n523), .Y(n383) );
  OAI21X1 U140 ( .A(n645), .B(n654), .C(n450), .Y(n384) );
  OAI21X1 U142 ( .A(n645), .B(n655), .C(n61), .Y(n385) );
  OAI21X1 U144 ( .A(n645), .B(n656), .C(n544), .Y(n386) );
  OAI21X1 U146 ( .A(n645), .B(n657), .C(n56), .Y(n387) );
  OAI21X1 U148 ( .A(n645), .B(n658), .C(n52), .Y(n388) );
  OAI21X1 U150 ( .A(n645), .B(n659), .C(n51), .Y(n389) );
  OAI21X1 U152 ( .A(n645), .B(n660), .C(n50), .Y(n390) );
  OAI21X1 U154 ( .A(n645), .B(n661), .C(n502), .Y(n391) );
  OAI21X1 U156 ( .A(n645), .B(n662), .C(n480), .Y(n392) );
  OAI21X1 U158 ( .A(n645), .B(n663), .C(n459), .Y(n393) );
  OAI21X1 U160 ( .A(n645), .B(n664), .C(n447), .Y(n394) );
  OAI21X1 U162 ( .A(n645), .B(n665), .C(n109), .Y(n395) );
  OAI21X1 U164 ( .A(n645), .B(n666), .C(n95), .Y(n396) );
  OAI21X1 U166 ( .A(n645), .B(n667), .C(n79), .Y(n397) );
  OAI21X1 U168 ( .A(n652), .B(n646), .C(n522), .Y(n398) );
  OAI21X1 U170 ( .A(n653), .B(n646), .C(n501), .Y(n399) );
  OAI21X1 U172 ( .A(n654), .B(n646), .C(n479), .Y(n400) );
  OAI21X1 U174 ( .A(n655), .B(n646), .C(n107), .Y(n401) );
  OAI21X1 U176 ( .A(n656), .B(n646), .C(n316), .Y(n402) );
  OAI21X1 U178 ( .A(n657), .B(n646), .C(n458), .Y(n403) );
  OAI21X1 U180 ( .A(n658), .B(n646), .C(n69), .Y(n404) );
  OAI21X1 U182 ( .A(n659), .B(n646), .C(n93), .Y(n405) );
  OAI21X1 U184 ( .A(n660), .B(n646), .C(n64), .Y(n406) );
  OAI21X1 U186 ( .A(n661), .B(n646), .C(n60), .Y(n407) );
  OAI21X1 U188 ( .A(n662), .B(n646), .C(n55), .Y(n408) );
  OAI21X1 U190 ( .A(n663), .B(n646), .C(n49), .Y(n409) );
  OAI21X1 U192 ( .A(n664), .B(n646), .C(n48), .Y(n410) );
  OAI21X1 U194 ( .A(n665), .B(n646), .C(n68), .Y(n411) );
  OAI21X1 U196 ( .A(n666), .B(n646), .C(n77), .Y(n412) );
  OAI21X1 U198 ( .A(n667), .B(n646), .C(n47), .Y(n413) );
  OAI21X1 U200 ( .A(n647), .B(n652), .C(n314), .Y(n414) );
  OAI21X1 U202 ( .A(n73), .B(n653), .C(n105), .Y(n415) );
  OAI21X1 U204 ( .A(n647), .B(n654), .C(n91), .Y(n416) );
  OAI21X1 U206 ( .A(n647), .B(n655), .C(n75), .Y(n417) );
  OAI21X1 U208 ( .A(n647), .B(n656), .C(n67), .Y(n418) );
  OAI21X1 U210 ( .A(n647), .B(n657), .C(n63), .Y(n419) );
  OAI21X1 U212 ( .A(n73), .B(n658), .C(n59), .Y(n420) );
  OAI21X1 U214 ( .A(n647), .B(n659), .C(n54), .Y(n421) );
  OAI21X1 U216 ( .A(n647), .B(n660), .C(n590), .Y(n422) );
  OAI21X1 U218 ( .A(n647), .B(n661), .C(n46), .Y(n423) );
  OAI21X1 U220 ( .A(n73), .B(n662), .C(n45), .Y(n424) );
  OAI21X1 U222 ( .A(n73), .B(n663), .C(n58), .Y(n425) );
  OAI21X1 U224 ( .A(n73), .B(n664), .C(n44), .Y(n426) );
  OAI21X1 U226 ( .A(n73), .B(n665), .C(n43), .Y(n427) );
  OAI21X1 U228 ( .A(n73), .B(n666), .C(n103), .Y(n428) );
  OAI21X1 U230 ( .A(n73), .B(n667), .C(n42), .Y(n429) );
  OAI21X1 U232 ( .A(n652), .B(n5), .C(n89), .Y(n430) );
  OAI21X1 U235 ( .A(n653), .B(n5), .C(n457), .Y(n431) );
  OAI21X1 U238 ( .A(n654), .B(n5), .C(n101), .Y(n432) );
  OAI21X1 U241 ( .A(n655), .B(n5), .C(n62), .Y(n433) );
  OAI21X1 U244 ( .A(n656), .B(n5), .C(n566), .Y(n434) );
  OAI21X1 U247 ( .A(n657), .B(n5), .C(n478), .Y(n435) );
  OAI21X1 U250 ( .A(n658), .B(n5), .C(n53), .Y(n436) );
  OAI21X1 U253 ( .A(n659), .B(n5), .C(n589), .Y(n437) );
  OAI21X1 U256 ( .A(n660), .B(n5), .C(n57), .Y(n438) );
  OAI21X1 U259 ( .A(n661), .B(n5), .C(n41), .Y(n439) );
  OAI21X1 U262 ( .A(n662), .B(n5), .C(n40), .Y(n440) );
  OAI21X1 U265 ( .A(n663), .B(n5), .C(n39), .Y(n441) );
  OAI21X1 U268 ( .A(n664), .B(n5), .C(n500), .Y(n442) );
  OAI21X1 U271 ( .A(n665), .B(n5), .C(n232), .Y(n443) );
  OAI21X1 U274 ( .A(n666), .B(n5), .C(n66), .Y(n444) );
  OAI21X1 U277 ( .A(n667), .B(n5), .C(n87), .Y(n445) );
  NAND3X1 U279 ( .A(n646), .B(n645), .C(n73), .Y(n143) );
  AOI22X1 U291 ( .A(n669), .B(r6[9]), .C(n672), .D(r7[9]), .Y(n228) );
  AOI22X1 U292 ( .A(n670), .B(r4[9]), .C(n673), .D(r5[9]), .Y(n227) );
  AOI22X1 U293 ( .A(n642), .B(r2[9]), .C(n644), .D(r3[9]), .Y(n225) );
  AOI22X1 U294 ( .A(n638), .B(r0[9]), .C(n640), .D(r1[9]), .Y(n224) );
  AOI22X1 U297 ( .A(n669), .B(r6[8]), .C(n672), .D(r7[8]), .Y(n241) );
  AOI22X1 U298 ( .A(n670), .B(r4[8]), .C(n673), .D(r5[8]), .Y(n240) );
  AOI22X1 U299 ( .A(n642), .B(r2[8]), .C(n644), .D(r3[8]), .Y(n238) );
  AOI22X1 U300 ( .A(n638), .B(r0[8]), .C(n640), .D(r1[8]), .Y(n237) );
  AOI22X1 U303 ( .A(n669), .B(r6[7]), .C(n672), .D(r7[7]), .Y(n246) );
  AOI22X1 U304 ( .A(n670), .B(r4[7]), .C(n673), .D(r5[7]), .Y(n245) );
  AOI22X1 U305 ( .A(n642), .B(r2[7]), .C(n644), .D(r3[7]), .Y(n243) );
  AOI22X1 U306 ( .A(n638), .B(r0[7]), .C(n640), .D(r1[7]), .Y(n242) );
  AOI22X1 U309 ( .A(n669), .B(r6[6]), .C(n672), .D(r7[6]), .Y(n251) );
  AOI22X1 U310 ( .A(n670), .B(r4[6]), .C(n673), .D(r5[6]), .Y(n250) );
  AOI22X1 U311 ( .A(n642), .B(r2[6]), .C(n644), .D(r3[6]), .Y(n248) );
  AOI22X1 U312 ( .A(n638), .B(r0[6]), .C(n640), .D(r1[6]), .Y(n247) );
  AOI22X1 U315 ( .A(n669), .B(r6[5]), .C(n672), .D(r7[5]), .Y(n256) );
  AOI22X1 U316 ( .A(n670), .B(r4[5]), .C(n673), .D(r5[5]), .Y(n255) );
  AOI22X1 U317 ( .A(n642), .B(r2[5]), .C(n644), .D(r3[5]), .Y(n253) );
  AOI22X1 U318 ( .A(n638), .B(r0[5]), .C(n640), .D(r1[5]), .Y(n252) );
  AOI22X1 U321 ( .A(n669), .B(r6[4]), .C(n672), .D(r7[4]), .Y(n261) );
  AOI22X1 U322 ( .A(n670), .B(r4[4]), .C(n673), .D(r5[4]), .Y(n260) );
  AOI22X1 U323 ( .A(n642), .B(r2[4]), .C(n644), .D(r3[4]), .Y(n258) );
  AOI22X1 U324 ( .A(n638), .B(r0[4]), .C(n640), .D(r1[4]), .Y(n257) );
  AOI22X1 U327 ( .A(n669), .B(r6[3]), .C(n672), .D(r7[3]), .Y(n266) );
  AOI22X1 U328 ( .A(n670), .B(r4[3]), .C(n673), .D(r5[3]), .Y(n265) );
  AOI22X1 U329 ( .A(n642), .B(r2[3]), .C(n644), .D(r3[3]), .Y(n263) );
  AOI22X1 U330 ( .A(n638), .B(r0[3]), .C(n640), .D(r1[3]), .Y(n262) );
  AOI22X1 U333 ( .A(n669), .B(r6[2]), .C(n672), .D(r7[2]), .Y(n271) );
  AOI22X1 U334 ( .A(n670), .B(r4[2]), .C(n673), .D(r5[2]), .Y(n270) );
  AOI22X1 U335 ( .A(n642), .B(r2[2]), .C(n644), .D(r3[2]), .Y(n268) );
  AOI22X1 U336 ( .A(n638), .B(r0[2]), .C(n640), .D(r1[2]), .Y(n267) );
  AOI22X1 U339 ( .A(n669), .B(r6[1]), .C(n672), .D(r7[1]), .Y(n276) );
  AOI22X1 U340 ( .A(n670), .B(r4[1]), .C(n673), .D(r5[1]), .Y(n275) );
  AOI22X1 U341 ( .A(n641), .B(r2[1]), .C(n643), .D(r3[1]), .Y(n273) );
  AOI22X1 U342 ( .A(n637), .B(r0[1]), .C(n639), .D(r1[1]), .Y(n272) );
  AOI22X1 U345 ( .A(n669), .B(r6[15]), .C(n672), .D(r7[15]), .Y(n281) );
  AOI22X1 U346 ( .A(n670), .B(r4[15]), .C(n673), .D(r5[15]), .Y(n280) );
  AOI22X1 U347 ( .A(n641), .B(r2[15]), .C(n643), .D(r3[15]), .Y(n278) );
  AOI22X1 U348 ( .A(n637), .B(r0[15]), .C(n639), .D(r1[15]), .Y(n277) );
  AOI22X1 U351 ( .A(n669), .B(r6[14]), .C(n672), .D(r7[14]), .Y(n286) );
  AOI22X1 U352 ( .A(n670), .B(r4[14]), .C(n673), .D(r5[14]), .Y(n285) );
  AOI22X1 U353 ( .A(n641), .B(r2[14]), .C(n643), .D(r3[14]), .Y(n283) );
  AOI22X1 U354 ( .A(n637), .B(r0[14]), .C(n639), .D(r1[14]), .Y(n282) );
  AOI22X1 U357 ( .A(n669), .B(r6[13]), .C(n672), .D(r7[13]), .Y(n291) );
  AOI22X1 U358 ( .A(n670), .B(r4[13]), .C(n673), .D(r5[13]), .Y(n290) );
  AOI22X1 U359 ( .A(n641), .B(r2[13]), .C(n643), .D(r3[13]), .Y(n288) );
  AOI22X1 U360 ( .A(n637), .B(r0[13]), .C(n639), .D(r1[13]), .Y(n287) );
  AOI22X1 U363 ( .A(n669), .B(r6[12]), .C(n672), .D(r7[12]), .Y(n296) );
  AOI22X1 U364 ( .A(n670), .B(r4[12]), .C(n673), .D(r5[12]), .Y(n295) );
  AOI22X1 U365 ( .A(n641), .B(r2[12]), .C(n643), .D(r3[12]), .Y(n293) );
  AOI22X1 U366 ( .A(n637), .B(r0[12]), .C(n639), .D(r1[12]), .Y(n292) );
  AOI22X1 U369 ( .A(n669), .B(r6[11]), .C(n672), .D(r7[11]), .Y(n301) );
  AOI22X1 U370 ( .A(n670), .B(r4[11]), .C(n673), .D(r5[11]), .Y(n300) );
  AOI22X1 U371 ( .A(n641), .B(r2[11]), .C(n643), .D(r3[11]), .Y(n298) );
  AOI22X1 U372 ( .A(n637), .B(r0[11]), .C(n639), .D(r1[11]), .Y(n297) );
  AOI22X1 U375 ( .A(n669), .B(r6[10]), .C(n672), .D(r7[10]), .Y(n306) );
  AOI22X1 U376 ( .A(n670), .B(r4[10]), .C(n673), .D(r5[10]), .Y(n305) );
  AOI22X1 U377 ( .A(n641), .B(r2[10]), .C(n643), .D(r3[10]), .Y(n303) );
  AOI22X1 U378 ( .A(n637), .B(r0[10]), .C(n639), .D(r1[10]), .Y(n302) );
  AOI22X1 U381 ( .A(n669), .B(r6[0]), .C(n672), .D(r7[0]), .Y(n311) );
  NAND3X1 U383 ( .A(readPtr[2]), .B(readPtr[1]), .C(readPtr[0]), .Y(n312) );
  NAND3X1 U385 ( .A(readPtr[1]), .B(n671), .C(readPtr[2]), .Y(n313) );
  AOI22X1 U386 ( .A(n670), .B(r4[0]), .C(n673), .D(r5[0]), .Y(n310) );
  NAND3X1 U388 ( .A(readPtr[2]), .B(n674), .C(readPtr[0]), .Y(n315) );
  NAND3X1 U390 ( .A(n671), .B(n674), .C(readPtr[2]), .Y(n317) );
  AOI22X1 U391 ( .A(n641), .B(r2[0]), .C(n643), .D(r3[0]), .Y(n308) );
  NOR3X1 U392 ( .A(n674), .B(readPtr[2]), .C(n671), .Y(n234) );
  NOR3X1 U393 ( .A(readPtr[0]), .B(readPtr[2]), .C(n674), .Y(n233) );
  AOI22X1 U395 ( .A(n637), .B(r0[0]), .C(n639), .D(r1[0]), .Y(n307) );
  NOR3X1 U396 ( .A(readPtr[1]), .B(readPtr[2]), .C(n671), .Y(n236) );
  NOR3X1 U398 ( .A(readPtr[1]), .B(readPtr[2]), .C(readPtr[0]), .Y(n235) );
  AND2X2 U400 ( .A(strobe[1]), .B(n599), .Y(n_0_net_) );
  AND2X1 U5 ( .A(n6), .B(n22), .Y(n309) );
  AND2X1 U7 ( .A(n13), .B(n29), .Y(n274) );
  AND2X1 U9 ( .A(n14), .B(n30), .Y(n269) );
  AND2X1 U11 ( .A(n15), .B(n31), .Y(n264) );
  AND2X1 U13 ( .A(n16), .B(n32), .Y(n259) );
  AND2X1 U15 ( .A(n17), .B(n33), .Y(n254) );
  AND2X1 U17 ( .A(n18), .B(n34), .Y(n249) );
  AND2X1 U19 ( .A(n19), .B(n35), .Y(n244) );
  AND2X1 U21 ( .A(n20), .B(n36), .Y(n239) );
  AND2X1 U23 ( .A(n21), .B(n37), .Y(n226) );
  AND2X1 U25 ( .A(n7), .B(n23), .Y(n304) );
  AND2X1 U27 ( .A(n8), .B(n24), .Y(n299) );
  AND2X1 U29 ( .A(n9), .B(n25), .Y(n294) );
  AND2X1 U31 ( .A(n10), .B(n26), .Y(n289) );
  AND2X1 U33 ( .A(n11), .B(n27), .Y(n284) );
  AND2X1 U35 ( .A(n12), .B(n28), .Y(n279) );
  AND2X1 U37 ( .A(n599), .B(n645), .Y(n448) );
  AND2X1 U39 ( .A(strobe[0]), .B(n599), .Y(n_1_net_) );
  OR2X1 U41 ( .A(n650), .B(n622), .Y(n73) );
  BUFX2 U43 ( .A(n317), .Y(n1) );
  BUFX2 U45 ( .A(n315), .Y(n2) );
  BUFX2 U47 ( .A(n313), .Y(n3) );
  BUFX2 U49 ( .A(n312), .Y(n4) );
  BUFX2 U51 ( .A(n143), .Y(n5) );
  OR2X1 U53 ( .A(n633), .B(n634), .Y(dout[8]) );
  OR2X1 U55 ( .A(n631), .B(n632), .Y(n634) );
  AND2X1 U57 ( .A(n574), .B(n622), .Y(n78) );
  AND2X1 U59 ( .A(n622), .B(n650), .Y(n76) );
  BUFX2 U61 ( .A(n310), .Y(n6) );
  BUFX2 U63 ( .A(n305), .Y(n7) );
  BUFX2 U65 ( .A(n300), .Y(n8) );
  BUFX2 U67 ( .A(n295), .Y(n9) );
  BUFX2 U69 ( .A(n290), .Y(n10) );
  BUFX2 U71 ( .A(n285), .Y(n11) );
  BUFX2 U73 ( .A(n280), .Y(n12) );
  BUFX2 U75 ( .A(n275), .Y(n13) );
  BUFX2 U77 ( .A(n270), .Y(n14) );
  BUFX2 U79 ( .A(n265), .Y(n15) );
  BUFX2 U81 ( .A(n260), .Y(n16) );
  BUFX2 U83 ( .A(n255), .Y(n17) );
  BUFX2 U85 ( .A(n250), .Y(n18) );
  BUFX2 U87 ( .A(n245), .Y(n19) );
  BUFX2 U89 ( .A(n240), .Y(n20) );
  BUFX2 U91 ( .A(n227), .Y(n21) );
  BUFX2 U93 ( .A(n311), .Y(n22) );
  BUFX2 U95 ( .A(n306), .Y(n23) );
  BUFX2 U97 ( .A(n301), .Y(n24) );
  BUFX2 U99 ( .A(n296), .Y(n25) );
  BUFX2 U101 ( .A(n291), .Y(n26) );
  BUFX2 U103 ( .A(n286), .Y(n27) );
  BUFX2 U105 ( .A(n281), .Y(n28) );
  BUFX2 U107 ( .A(n276), .Y(n29) );
  BUFX2 U109 ( .A(n271), .Y(n30) );
  BUFX2 U111 ( .A(n266), .Y(n31) );
  BUFX2 U113 ( .A(n261), .Y(n32) );
  BUFX2 U115 ( .A(n256), .Y(n33) );
  BUFX2 U117 ( .A(n251), .Y(n34) );
  BUFX2 U119 ( .A(n246), .Y(n35) );
  BUFX2 U121 ( .A(n241), .Y(n36) );
  BUFX2 U123 ( .A(n228), .Y(n37) );
  BUFX2 U125 ( .A(n74), .Y(n38) );
  AND2X1 U127 ( .A(r0[11]), .B(n5), .Y(n219) );
  INVX1 U129 ( .A(n219), .Y(n39) );
  AND2X1 U131 ( .A(r0[10]), .B(n5), .Y(n218) );
  INVX1 U133 ( .A(n218), .Y(n40) );
  AND2X1 U135 ( .A(r0[9]), .B(n5), .Y(n217) );
  INVX1 U137 ( .A(n217), .Y(n41) );
  AND2X1 U139 ( .A(r2[15]), .B(n647), .Y(n207) );
  INVX1 U141 ( .A(n207), .Y(n42) );
  AND2X1 U143 ( .A(r2[13]), .B(n647), .Y(n205) );
  INVX1 U145 ( .A(n205), .Y(n43) );
  AND2X1 U147 ( .A(r2[12]), .B(n647), .Y(n204) );
  INVX1 U149 ( .A(n204), .Y(n44) );
  AND2X1 U151 ( .A(r2[10]), .B(n647), .Y(n202) );
  INVX1 U153 ( .A(n202), .Y(n45) );
  AND2X1 U155 ( .A(r2[9]), .B(n647), .Y(n201) );
  INVX1 U157 ( .A(n201), .Y(n46) );
  AND2X1 U159 ( .A(r4[15]), .B(n646), .Y(n191) );
  INVX1 U161 ( .A(n191), .Y(n47) );
  AND2X1 U163 ( .A(r4[12]), .B(n646), .Y(n188) );
  INVX1 U165 ( .A(n188), .Y(n48) );
  AND2X1 U167 ( .A(r4[11]), .B(n646), .Y(n187) );
  INVX1 U169 ( .A(n187), .Y(n49) );
  AND2X1 U171 ( .A(r6[8]), .B(n645), .Y(n168) );
  INVX1 U173 ( .A(n168), .Y(n50) );
  AND2X1 U175 ( .A(r6[7]), .B(n645), .Y(n167) );
  INVX1 U177 ( .A(n167), .Y(n51) );
  AND2X1 U179 ( .A(r6[6]), .B(n645), .Y(n166) );
  INVX1 U181 ( .A(n166), .Y(n52) );
  OR2X1 U183 ( .A(n511), .B(n512), .Y(dout[15]) );
  OR2X1 U185 ( .A(n509), .B(n510), .Y(n512) );
  AND2X1 U187 ( .A(r0[6]), .B(n5), .Y(n214) );
  INVX1 U189 ( .A(n214), .Y(n53) );
  AND2X1 U191 ( .A(r2[7]), .B(n647), .Y(n199) );
  INVX1 U193 ( .A(n199), .Y(n54) );
  AND2X1 U195 ( .A(r4[10]), .B(n646), .Y(n186) );
  INVX1 U197 ( .A(n186), .Y(n55) );
  AND2X1 U199 ( .A(r6[5]), .B(n645), .Y(n165) );
  INVX1 U201 ( .A(n165), .Y(n56) );
  OR2X1 U203 ( .A(n474), .B(n475), .Y(dout[7]) );
  OR2X1 U205 ( .A(n472), .B(n473), .Y(n475) );
  OR2X1 U207 ( .A(n562), .B(n563), .Y(dout[10]) );
  OR2X1 U209 ( .A(n560), .B(n561), .Y(n563) );
  AND2X1 U211 ( .A(r0[8]), .B(n5), .Y(n216) );
  INVX1 U213 ( .A(n216), .Y(n57) );
  AND2X1 U215 ( .A(r2[11]), .B(n647), .Y(n203) );
  INVX1 U217 ( .A(n203), .Y(n58) );
  AND2X1 U219 ( .A(r2[6]), .B(n647), .Y(n198) );
  INVX1 U221 ( .A(n198), .Y(n59) );
  AND2X1 U223 ( .A(r4[9]), .B(n646), .Y(n185) );
  INVX1 U225 ( .A(n185), .Y(n60) );
  AND2X1 U227 ( .A(r6[3]), .B(n645), .Y(n163) );
  INVX1 U229 ( .A(n163), .Y(n61) );
  OR2X1 U231 ( .A(n518), .B(n519), .Y(dout[2]) );
  OR2X1 U233 ( .A(n516), .B(n517), .Y(n519) );
  OR2X1 U234 ( .A(n610), .B(n611), .Y(dout[12]) );
  OR2X1 U236 ( .A(n608), .B(n609), .Y(n611) );
  AND2X1 U237 ( .A(r0[3]), .B(n5), .Y(n211) );
  INVX1 U239 ( .A(n211), .Y(n62) );
  AND2X1 U240 ( .A(r2[5]), .B(n647), .Y(n197) );
  INVX1 U242 ( .A(n197), .Y(n63) );
  AND2X1 U243 ( .A(r4[8]), .B(n646), .Y(n184) );
  INVX1 U245 ( .A(n184), .Y(n64) );
  AND2X1 U246 ( .A(r6[0]), .B(n645), .Y(n160) );
  INVX1 U248 ( .A(n160), .Y(n65) );
  OR2X1 U249 ( .A(n540), .B(n541), .Y(dout[3]) );
  OR2X1 U251 ( .A(n538), .B(n539), .Y(n541) );
  OR2X1 U252 ( .A(n585), .B(n586), .Y(dout[11]) );
  OR2X1 U254 ( .A(n583), .B(n584), .Y(n586) );
  AND2X1 U255 ( .A(r0[14]), .B(n5), .Y(n222) );
  INVX1 U257 ( .A(n222), .Y(n66) );
  AND2X1 U258 ( .A(r2[4]), .B(n647), .Y(n196) );
  INVX1 U260 ( .A(n196), .Y(n67) );
  AND2X1 U261 ( .A(r4[13]), .B(n646), .Y(n189) );
  INVX1 U263 ( .A(n189), .Y(n68) );
  AND2X1 U264 ( .A(r4[6]), .B(n646), .Y(n182) );
  INVX1 U266 ( .A(n182), .Y(n69) );
  AND2X1 U267 ( .A(r1[12]), .B(n5), .Y(n156) );
  INVX1 U269 ( .A(n156), .Y(n70) );
  AND2X1 U270 ( .A(r7[15]), .B(n645), .Y(n110) );
  INVX1 U272 ( .A(n110), .Y(n71) );
  OR2X1 U273 ( .A(n555), .B(n556), .Y(dout[4]) );
  OR2X1 U275 ( .A(n553), .B(n554), .Y(n556) );
  OR2X1 U276 ( .A(n626), .B(n627), .Y(dout[13]) );
  OR2X1 U278 ( .A(n624), .B(n625), .Y(n627) );
  AND2X1 U280 ( .A(r2[3]), .B(n647), .Y(n195) );
  INVX1 U281 ( .A(n195), .Y(n75) );
  AND2X1 U282 ( .A(r4[14]), .B(n646), .Y(n190) );
  INVX1 U283 ( .A(n190), .Y(n77) );
  AND2X1 U284 ( .A(r6[15]), .B(n645), .Y(n175) );
  INVX1 U285 ( .A(n175), .Y(n79) );
  AND2X1 U286 ( .A(r1[11]), .B(n5), .Y(n155) );
  INVX1 U287 ( .A(n155), .Y(n81) );
  AND2X1 U288 ( .A(r5[12]), .B(n646), .Y(n123) );
  INVX1 U289 ( .A(n123), .Y(n83) );
  AND2X1 U290 ( .A(r7[13]), .B(n645), .Y(n106) );
  INVX1 U295 ( .A(n106), .Y(n85) );
  OR2X1 U296 ( .A(n578), .B(n579), .Y(dout[5]) );
  OR2X1 U301 ( .A(n576), .B(n577), .Y(n579) );
  OR2X1 U302 ( .A(n533), .B(n534), .Y(dout[14]) );
  OR2X1 U307 ( .A(n531), .B(n532), .Y(n534) );
  AND2X1 U308 ( .A(r0[15]), .B(n5), .Y(n223) );
  INVX1 U313 ( .A(n223), .Y(n87) );
  AND2X1 U314 ( .A(r0[0]), .B(n5), .Y(n208) );
  INVX1 U319 ( .A(n208), .Y(n89) );
  AND2X1 U320 ( .A(r2[2]), .B(n647), .Y(n194) );
  INVX1 U325 ( .A(n194), .Y(n91) );
  AND2X1 U326 ( .A(r4[7]), .B(n646), .Y(n183) );
  INVX1 U331 ( .A(n183), .Y(n93) );
  AND2X1 U332 ( .A(r6[14]), .B(n645), .Y(n174) );
  INVX1 U337 ( .A(n174), .Y(n95) );
  AND2X1 U338 ( .A(r5[11]), .B(n646), .Y(n122) );
  INVX1 U343 ( .A(n122), .Y(n97) );
  AND2X1 U344 ( .A(r7[12]), .B(n645), .Y(n104) );
  INVX1 U349 ( .A(n104), .Y(n99) );
  OR2X1 U350 ( .A(n496), .B(n497), .Y(dout[6]) );
  OR2X1 U355 ( .A(n494), .B(n495), .Y(n497) );
  OR2X1 U356 ( .A(n467), .B(n468), .Y(dout[0]) );
  OR2X1 U361 ( .A(n465), .B(n466), .Y(n468) );
  AND2X1 U362 ( .A(r0[2]), .B(n5), .Y(n210) );
  INVX1 U367 ( .A(n210), .Y(n101) );
  AND2X1 U368 ( .A(r2[14]), .B(n647), .Y(n206) );
  INVX1 U373 ( .A(n206), .Y(n103) );
  AND2X1 U374 ( .A(r2[1]), .B(n647), .Y(n193) );
  INVX1 U379 ( .A(n193), .Y(n105) );
  AND2X1 U380 ( .A(r4[3]), .B(n646), .Y(n179) );
  INVX1 U382 ( .A(n179), .Y(n107) );
  AND2X1 U384 ( .A(r6[13]), .B(n645), .Y(n173) );
  INVX1 U387 ( .A(n173), .Y(n109) );
  AND2X1 U389 ( .A(r1[10]), .B(n5), .Y(n154) );
  INVX1 U394 ( .A(n154), .Y(n229) );
  AND2X1 U397 ( .A(r5[9]), .B(n646), .Y(n120) );
  INVX1 U399 ( .A(n120), .Y(n230) );
  AND2X1 U403 ( .A(r7[11]), .B(n645), .Y(n102) );
  INVX1 U404 ( .A(n102), .Y(n231) );
  OR2X1 U405 ( .A(n603), .B(n604), .Y(dout[9]) );
  OR2X1 U406 ( .A(n601), .B(n602), .Y(n604) );
  OR2X1 U407 ( .A(n489), .B(n490), .Y(dout[1]) );
  OR2X1 U408 ( .A(n487), .B(n488), .Y(n490) );
  AND2X1 U409 ( .A(r0[13]), .B(n5), .Y(n221) );
  INVX1 U410 ( .A(n221), .Y(n232) );
  AND2X1 U411 ( .A(r2[0]), .B(n647), .Y(n192) );
  INVX1 U412 ( .A(n192), .Y(n314) );
  AND2X1 U413 ( .A(r4[4]), .B(n646), .Y(n180) );
  INVX1 U414 ( .A(n180), .Y(n316) );
  AND2X1 U415 ( .A(r6[12]), .B(n645), .Y(n172) );
  INVX1 U416 ( .A(n172), .Y(n447) );
  AND2X1 U417 ( .A(r6[2]), .B(n645), .Y(n162) );
  INVX1 U418 ( .A(n162), .Y(n450) );
  AND2X1 U419 ( .A(r1[6]), .B(n5), .Y(n150) );
  INVX1 U420 ( .A(n150), .Y(n451) );
  AND2X1 U421 ( .A(r3[8]), .B(n73), .Y(n135) );
  INVX1 U422 ( .A(n135), .Y(n454) );
  AND2X1 U423 ( .A(r5[10]), .B(n646), .Y(n121) );
  INVX1 U424 ( .A(n121), .Y(n455) );
  AND2X1 U425 ( .A(r7[9]), .B(n645), .Y(n98) );
  INVX1 U426 ( .A(n98), .Y(n456) );
  AND2X1 U427 ( .A(r0[1]), .B(n5), .Y(n209) );
  INVX1 U428 ( .A(n209), .Y(n457) );
  AND2X1 U429 ( .A(r4[5]), .B(n646), .Y(n181) );
  INVX1 U430 ( .A(n181), .Y(n458) );
  AND2X1 U431 ( .A(r6[11]), .B(n645), .Y(n171) );
  INVX1 U432 ( .A(n171), .Y(n459) );
  AND2X1 U433 ( .A(r1[4]), .B(n5), .Y(n148) );
  INVX1 U434 ( .A(n148), .Y(n460) );
  AND2X1 U435 ( .A(r3[15]), .B(n647), .Y(n142) );
  INVX1 U436 ( .A(n142), .Y(n461) );
  AND2X1 U437 ( .A(r5[7]), .B(n646), .Y(n118) );
  INVX1 U438 ( .A(n118), .Y(n462) );
  AND2X1 U439 ( .A(r7[8]), .B(n645), .Y(n96) );
  INVX1 U440 ( .A(n96), .Y(n463) );
  INVX1 U441 ( .A(n309), .Y(n465) );
  INVX1 U442 ( .A(n470), .Y(n466) );
  INVX1 U443 ( .A(n469), .Y(n467) );
  BUFX2 U444 ( .A(n307), .Y(n469) );
  BUFX2 U445 ( .A(n308), .Y(n470) );
  INVX1 U446 ( .A(n244), .Y(n472) );
  INVX1 U447 ( .A(n477), .Y(n473) );
  INVX1 U448 ( .A(n476), .Y(n474) );
  BUFX2 U449 ( .A(n242), .Y(n476) );
  BUFX2 U450 ( .A(n243), .Y(n477) );
  AND2X1 U451 ( .A(r0[5]), .B(n5), .Y(n213) );
  INVX1 U452 ( .A(n213), .Y(n478) );
  AND2X1 U453 ( .A(r4[2]), .B(n646), .Y(n178) );
  INVX1 U454 ( .A(n178), .Y(n479) );
  AND2X1 U455 ( .A(r6[10]), .B(n645), .Y(n170) );
  INVX1 U456 ( .A(n170), .Y(n480) );
  AND2X1 U457 ( .A(r1[9]), .B(n5), .Y(n153) );
  INVX1 U458 ( .A(n153), .Y(n481) );
  AND2X1 U459 ( .A(r3[14]), .B(n647), .Y(n141) );
  INVX1 U460 ( .A(n141), .Y(n482) );
  AND2X1 U461 ( .A(r3[4]), .B(n647), .Y(n131) );
  INVX1 U462 ( .A(n131), .Y(n483) );
  AND2X1 U463 ( .A(r5[8]), .B(n646), .Y(n119) );
  INVX1 U464 ( .A(n119), .Y(n484) );
  AND2X1 U465 ( .A(r7[7]), .B(n645), .Y(n94) );
  INVX1 U466 ( .A(n94), .Y(n485) );
  INVX1 U467 ( .A(n274), .Y(n487) );
  INVX1 U468 ( .A(n492), .Y(n488) );
  INVX1 U469 ( .A(n491), .Y(n489) );
  BUFX2 U470 ( .A(n272), .Y(n491) );
  BUFX2 U471 ( .A(n273), .Y(n492) );
  INVX1 U472 ( .A(n249), .Y(n494) );
  INVX1 U473 ( .A(n499), .Y(n495) );
  INVX1 U474 ( .A(n498), .Y(n496) );
  BUFX2 U475 ( .A(n247), .Y(n498) );
  BUFX2 U476 ( .A(n248), .Y(n499) );
  AND2X1 U477 ( .A(r0[12]), .B(n5), .Y(n220) );
  INVX1 U478 ( .A(n220), .Y(n500) );
  AND2X1 U479 ( .A(r4[1]), .B(n646), .Y(n177) );
  INVX1 U480 ( .A(n177), .Y(n501) );
  AND2X1 U481 ( .A(r6[9]), .B(n645), .Y(n169) );
  INVX1 U482 ( .A(n169), .Y(n502) );
  AND2X1 U483 ( .A(r1[8]), .B(n5), .Y(n152) );
  INVX1 U484 ( .A(n152), .Y(n503) );
  AND2X1 U485 ( .A(r3[13]), .B(n647), .Y(n140) );
  INVX1 U486 ( .A(n140), .Y(n504) );
  AND2X1 U487 ( .A(r3[5]), .B(n647), .Y(n132) );
  INVX1 U488 ( .A(n132), .Y(n505) );
  AND2X1 U489 ( .A(r5[4]), .B(n646), .Y(n115) );
  INVX1 U490 ( .A(n115), .Y(n506) );
  AND2X1 U491 ( .A(r7[6]), .B(n645), .Y(n92) );
  INVX1 U492 ( .A(n92), .Y(n507) );
  INVX1 U493 ( .A(n279), .Y(n509) );
  INVX1 U494 ( .A(n514), .Y(n510) );
  INVX1 U495 ( .A(n513), .Y(n511) );
  BUFX2 U496 ( .A(n277), .Y(n513) );
  BUFX2 U497 ( .A(n278), .Y(n514) );
  INVX1 U498 ( .A(n269), .Y(n516) );
  INVX1 U499 ( .A(n521), .Y(n517) );
  INVX1 U500 ( .A(n520), .Y(n518) );
  BUFX2 U501 ( .A(n267), .Y(n520) );
  BUFX2 U502 ( .A(n268), .Y(n521) );
  AND2X1 U503 ( .A(r4[0]), .B(n646), .Y(n176) );
  INVX1 U504 ( .A(n176), .Y(n522) );
  AND2X1 U505 ( .A(r6[1]), .B(n645), .Y(n161) );
  INVX1 U506 ( .A(n161), .Y(n523) );
  AND2X1 U507 ( .A(r1[15]), .B(n5), .Y(n159) );
  INVX1 U508 ( .A(n159), .Y(n524) );
  AND2X1 U509 ( .A(r1[7]), .B(n5), .Y(n151) );
  INVX1 U510 ( .A(n151), .Y(n525) );
  AND2X1 U511 ( .A(r3[10]), .B(n647), .Y(n137) );
  INVX1 U512 ( .A(n137), .Y(n526) );
  AND2X1 U513 ( .A(r3[6]), .B(n73), .Y(n133) );
  INVX1 U514 ( .A(n133), .Y(n527) );
  AND2X1 U515 ( .A(r5[5]), .B(n646), .Y(n116) );
  INVX1 U516 ( .A(n116), .Y(n528) );
  AND2X1 U517 ( .A(r7[4]), .B(n645), .Y(n88) );
  INVX1 U518 ( .A(n88), .Y(n529) );
  INVX1 U519 ( .A(n284), .Y(n531) );
  INVX1 U520 ( .A(n536), .Y(n532) );
  INVX1 U521 ( .A(n535), .Y(n533) );
  BUFX2 U522 ( .A(n282), .Y(n535) );
  BUFX2 U523 ( .A(n283), .Y(n536) );
  INVX1 U524 ( .A(n264), .Y(n538) );
  INVX1 U525 ( .A(n543), .Y(n539) );
  INVX1 U526 ( .A(n542), .Y(n540) );
  BUFX2 U527 ( .A(n262), .Y(n542) );
  BUFX2 U528 ( .A(n263), .Y(n543) );
  AND2X1 U529 ( .A(r6[4]), .B(n645), .Y(n164) );
  INVX1 U530 ( .A(n164), .Y(n544) );
  AND2X1 U531 ( .A(r1[5]), .B(n5), .Y(n149) );
  INVX1 U532 ( .A(n149), .Y(n545) );
  AND2X1 U533 ( .A(r1[0]), .B(n5), .Y(n144) );
  INVX1 U534 ( .A(n144), .Y(n546) );
  AND2X1 U535 ( .A(r3[12]), .B(n647), .Y(n139) );
  INVX1 U536 ( .A(n139), .Y(n547) );
  AND2X1 U537 ( .A(r3[1]), .B(n647), .Y(n128) );
  INVX1 U538 ( .A(n128), .Y(n548) );
  AND2X1 U539 ( .A(r5[14]), .B(n646), .Y(n125) );
  INVX1 U540 ( .A(n125), .Y(n549) );
  AND2X1 U541 ( .A(r5[2]), .B(n646), .Y(n113) );
  INVX1 U542 ( .A(n113), .Y(n550) );
  AND2X1 U543 ( .A(r7[3]), .B(n645), .Y(n86) );
  INVX1 U544 ( .A(n86), .Y(n551) );
  INVX1 U545 ( .A(n259), .Y(n553) );
  INVX1 U546 ( .A(n558), .Y(n554) );
  INVX1 U547 ( .A(n557), .Y(n555) );
  BUFX2 U548 ( .A(n257), .Y(n557) );
  BUFX2 U549 ( .A(n258), .Y(n558) );
  INVX1 U550 ( .A(n304), .Y(n560) );
  INVX1 U551 ( .A(n565), .Y(n561) );
  INVX1 U552 ( .A(n564), .Y(n562) );
  BUFX2 U553 ( .A(n302), .Y(n564) );
  BUFX2 U554 ( .A(n303), .Y(n565) );
  AND2X1 U555 ( .A(r0[4]), .B(n5), .Y(n212) );
  INVX1 U556 ( .A(n212), .Y(n566) );
  AND2X1 U557 ( .A(r1[1]), .B(n5), .Y(n145) );
  INVX1 U558 ( .A(n145), .Y(n567) );
  AND2X1 U559 ( .A(r3[9]), .B(n647), .Y(n136) );
  INVX1 U560 ( .A(n136), .Y(n568) );
  AND2X1 U561 ( .A(r3[0]), .B(n647), .Y(n127) );
  INVX1 U562 ( .A(n127), .Y(n569) );
  AND2X1 U563 ( .A(r5[15]), .B(n646), .Y(n126) );
  INVX1 U564 ( .A(n126), .Y(n570) );
  AND2X1 U565 ( .A(r5[3]), .B(n646), .Y(n114) );
  INVX1 U566 ( .A(n114), .Y(n571) );
  AND2X1 U567 ( .A(r7[14]), .B(n645), .Y(n108) );
  INVX1 U568 ( .A(n108), .Y(n572) );
  AND2X1 U569 ( .A(r7[2]), .B(n645), .Y(n84) );
  INVX1 U570 ( .A(n84), .Y(n573) );
  BUFX2 U571 ( .A(count[0]), .Y(n574) );
  INVX1 U572 ( .A(n254), .Y(n576) );
  INVX1 U573 ( .A(n581), .Y(n577) );
  INVX1 U574 ( .A(n580), .Y(n578) );
  BUFX2 U575 ( .A(n252), .Y(n580) );
  BUFX2 U576 ( .A(n253), .Y(n581) );
  INVX1 U577 ( .A(n299), .Y(n583) );
  INVX1 U578 ( .A(n588), .Y(n584) );
  INVX1 U579 ( .A(n587), .Y(n585) );
  BUFX2 U580 ( .A(n297), .Y(n587) );
  BUFX2 U581 ( .A(n298), .Y(n588) );
  AND2X1 U582 ( .A(r0[7]), .B(n5), .Y(n215) );
  INVX1 U583 ( .A(n215), .Y(n589) );
  AND2X1 U584 ( .A(r2[8]), .B(n647), .Y(n200) );
  INVX1 U585 ( .A(n200), .Y(n590) );
  AND2X1 U586 ( .A(r1[13]), .B(n5), .Y(n157) );
  INVX1 U587 ( .A(n157), .Y(n591) );
  AND2X1 U588 ( .A(r1[2]), .B(n5), .Y(n146) );
  INVX1 U589 ( .A(n146), .Y(n592) );
  AND2X1 U590 ( .A(r3[11]), .B(n647), .Y(n138) );
  INVX1 U591 ( .A(n138), .Y(n593) );
  AND2X1 U592 ( .A(r3[3]), .B(n647), .Y(n130) );
  INVX1 U593 ( .A(n130), .Y(n594) );
  AND2X1 U594 ( .A(r5[6]), .B(n646), .Y(n117) );
  INVX1 U595 ( .A(n117), .Y(n595) );
  AND2X1 U596 ( .A(r5[0]), .B(n646), .Y(n111) );
  INVX1 U597 ( .A(n111), .Y(n596) );
  AND2X1 U598 ( .A(r7[10]), .B(n645), .Y(n100) );
  INVX1 U599 ( .A(n100), .Y(n597) );
  AND2X1 U600 ( .A(r7[1]), .B(n645), .Y(n82) );
  INVX1 U601 ( .A(n82), .Y(n598) );
  BUFX2 U602 ( .A(F0), .Y(n599) );
  INVX1 U603 ( .A(n226), .Y(n601) );
  INVX1 U604 ( .A(n606), .Y(n602) );
  INVX1 U605 ( .A(n605), .Y(n603) );
  BUFX2 U606 ( .A(n224), .Y(n605) );
  BUFX2 U607 ( .A(n225), .Y(n606) );
  INVX1 U608 ( .A(n294), .Y(n608) );
  INVX1 U609 ( .A(n613), .Y(n609) );
  INVX1 U610 ( .A(n612), .Y(n610) );
  BUFX2 U611 ( .A(n292), .Y(n612) );
  BUFX2 U612 ( .A(n293), .Y(n613) );
  AND2X1 U613 ( .A(r1[14]), .B(n5), .Y(n158) );
  INVX1 U614 ( .A(n158), .Y(n614) );
  AND2X1 U615 ( .A(r1[3]), .B(n5), .Y(n147) );
  INVX1 U616 ( .A(n147), .Y(n615) );
  AND2X1 U617 ( .A(r3[7]), .B(n647), .Y(n134) );
  INVX1 U618 ( .A(n134), .Y(n616) );
  AND2X1 U619 ( .A(r3[2]), .B(n73), .Y(n129) );
  INVX1 U620 ( .A(n129), .Y(n617) );
  AND2X1 U621 ( .A(r5[13]), .B(n646), .Y(n124) );
  INVX1 U622 ( .A(n124), .Y(n618) );
  AND2X1 U623 ( .A(r5[1]), .B(n646), .Y(n112) );
  INVX1 U624 ( .A(n112), .Y(n619) );
  AND2X1 U625 ( .A(r7[5]), .B(n645), .Y(n90) );
  INVX1 U626 ( .A(n90), .Y(n620) );
  AND2X1 U627 ( .A(r7[0]), .B(n645), .Y(n80) );
  INVX1 U628 ( .A(n80), .Y(n621) );
  BUFX2 U629 ( .A(count[1]), .Y(n622) );
  INVX1 U630 ( .A(n289), .Y(n624) );
  INVX1 U631 ( .A(n629), .Y(n625) );
  INVX1 U632 ( .A(n628), .Y(n626) );
  BUFX2 U633 ( .A(n287), .Y(n628) );
  BUFX2 U634 ( .A(n288), .Y(n629) );
  INVX1 U635 ( .A(n239), .Y(n631) );
  INVX1 U636 ( .A(n636), .Y(n632) );
  INVX1 U637 ( .A(n635), .Y(n633) );
  BUFX2 U638 ( .A(n237), .Y(n635) );
  BUFX2 U639 ( .A(n238), .Y(n636) );
  INVX1 U640 ( .A(reset), .Y(n649) );
  INVX1 U641 ( .A(n648), .Y(n647) );
  INVX1 U642 ( .A(n78), .Y(n645) );
  INVX1 U643 ( .A(n76), .Y(n646) );
  BUFX2 U644 ( .A(n234), .Y(n643) );
  BUFX2 U645 ( .A(n234), .Y(n644) );
  BUFX2 U646 ( .A(n236), .Y(n639) );
  BUFX2 U647 ( .A(n236), .Y(n640) );
  BUFX2 U648 ( .A(n233), .Y(n641) );
  BUFX2 U649 ( .A(n233), .Y(n642) );
  BUFX2 U650 ( .A(n235), .Y(n637) );
  BUFX2 U651 ( .A(n235), .Y(n638) );
  INVX1 U652 ( .A(n73), .Y(n648) );
  AND2X1 U653 ( .A(listen), .B(n649), .Y(n72) );
  INVX1 U654 ( .A(din[0]), .Y(n652) );
  INVX1 U655 ( .A(din[1]), .Y(n653) );
  INVX1 U656 ( .A(din[2]), .Y(n654) );
  INVX1 U657 ( .A(din[3]), .Y(n655) );
  INVX1 U658 ( .A(din[4]), .Y(n656) );
  INVX1 U659 ( .A(din[5]), .Y(n657) );
  INVX1 U660 ( .A(din[6]), .Y(n658) );
  INVX1 U661 ( .A(din[7]), .Y(n659) );
  INVX1 U662 ( .A(din[8]), .Y(n660) );
  INVX1 U663 ( .A(din[9]), .Y(n661) );
  INVX1 U664 ( .A(din[10]), .Y(n662) );
  INVX1 U665 ( .A(din[11]), .Y(n663) );
  INVX1 U666 ( .A(din[12]), .Y(n664) );
  INVX1 U667 ( .A(din[13]), .Y(n665) );
  INVX1 U668 ( .A(din[14]), .Y(n666) );
  INVX1 U669 ( .A(din[15]), .Y(n667) );
  INVX1 U670 ( .A(n2), .Y(n673) );
  INVX1 U671 ( .A(n4), .Y(n672) );
  INVX1 U672 ( .A(n3), .Y(n669) );
  INVX1 U673 ( .A(n1), .Y(n670) );
  INVX1 U674 ( .A(readPtr[1]), .Y(n674) );
  INVX1 U675 ( .A(readPtr[0]), .Y(n671) );
  INVX1 U676 ( .A(n574), .Y(n650) );
  INVX1 U677 ( .A(listen), .Y(n668) );
  INVX1 U678 ( .A(dStrobe0), .Y(n651) );
endmodule


module Processing_logic_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [15:1] carry;

  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YC(carry[15]), .YS(
        SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(carry[1]), .YC(carry[2]), .YS(SUM[1]) );
  AND2X1 U1 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
  XOR2X1 U2 ( .A(B[15]), .B(A[15]), .Y(n1) );
  XOR2X1 U3 ( .A(carry[15]), .B(n1), .Y(SUM[15]) );
  XOR2X1 U4 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module Processing_logic_DW01_add_2 ( A, B, CI, SUM, CO );
  input [25:0] A;
  input [25:0] B;
  output [25:0] SUM;
  input CI;
  output CO;

  wire   [25:5] carry;
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign SUM[0] = A[0];

  INVX1 U1 ( .A(A[3]), .Y(SUM[3]) );
  XOR2X1 U2 ( .A(A[25]), .B(carry[25]), .Y(SUM[25]) );
  AND2X1 U3 ( .A(carry[24]), .B(A[24]), .Y(carry[25]) );
  XOR2X1 U4 ( .A(carry[24]), .B(A[24]), .Y(SUM[24]) );
  AND2X1 U5 ( .A(carry[23]), .B(A[23]), .Y(carry[24]) );
  XOR2X1 U6 ( .A(carry[23]), .B(A[23]), .Y(SUM[23]) );
  AND2X1 U7 ( .A(carry[22]), .B(A[22]), .Y(carry[23]) );
  XOR2X1 U8 ( .A(carry[22]), .B(A[22]), .Y(SUM[22]) );
  AND2X1 U9 ( .A(carry[21]), .B(A[21]), .Y(carry[22]) );
  XOR2X1 U10 ( .A(carry[21]), .B(A[21]), .Y(SUM[21]) );
  AND2X1 U11 ( .A(carry[20]), .B(A[20]), .Y(carry[21]) );
  XOR2X1 U12 ( .A(carry[20]), .B(A[20]), .Y(SUM[20]) );
  AND2X1 U13 ( .A(carry[19]), .B(A[19]), .Y(carry[20]) );
  XOR2X1 U14 ( .A(carry[19]), .B(A[19]), .Y(SUM[19]) );
  AND2X1 U15 ( .A(carry[18]), .B(A[18]), .Y(carry[19]) );
  XOR2X1 U16 ( .A(carry[18]), .B(A[18]), .Y(SUM[18]) );
  AND2X1 U17 ( .A(carry[17]), .B(A[17]), .Y(carry[18]) );
  XOR2X1 U18 ( .A(carry[17]), .B(A[17]), .Y(SUM[17]) );
  AND2X1 U19 ( .A(carry[16]), .B(A[16]), .Y(carry[17]) );
  XOR2X1 U20 ( .A(carry[16]), .B(A[16]), .Y(SUM[16]) );
  AND2X1 U21 ( .A(carry[15]), .B(A[15]), .Y(carry[16]) );
  XOR2X1 U22 ( .A(carry[15]), .B(A[15]), .Y(SUM[15]) );
  AND2X1 U23 ( .A(carry[14]), .B(A[14]), .Y(carry[15]) );
  XOR2X1 U24 ( .A(carry[14]), .B(A[14]), .Y(SUM[14]) );
  AND2X1 U25 ( .A(carry[13]), .B(A[13]), .Y(carry[14]) );
  XOR2X1 U26 ( .A(carry[13]), .B(A[13]), .Y(SUM[13]) );
  AND2X1 U27 ( .A(carry[12]), .B(A[12]), .Y(carry[13]) );
  XOR2X1 U28 ( .A(carry[12]), .B(A[12]), .Y(SUM[12]) );
  AND2X1 U29 ( .A(carry[11]), .B(A[11]), .Y(carry[12]) );
  XOR2X1 U30 ( .A(carry[11]), .B(A[11]), .Y(SUM[11]) );
  AND2X1 U31 ( .A(carry[10]), .B(A[10]), .Y(carry[11]) );
  XOR2X1 U32 ( .A(carry[10]), .B(A[10]), .Y(SUM[10]) );
  AND2X1 U33 ( .A(carry[9]), .B(A[9]), .Y(carry[10]) );
  XOR2X1 U34 ( .A(carry[9]), .B(A[9]), .Y(SUM[9]) );
  AND2X1 U35 ( .A(carry[8]), .B(A[8]), .Y(carry[9]) );
  XOR2X1 U36 ( .A(carry[8]), .B(A[8]), .Y(SUM[8]) );
  AND2X1 U37 ( .A(carry[7]), .B(A[7]), .Y(carry[8]) );
  XOR2X1 U38 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  AND2X1 U39 ( .A(carry[6]), .B(A[6]), .Y(carry[7]) );
  XOR2X1 U40 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  AND2X1 U41 ( .A(carry[5]), .B(A[5]), .Y(carry[6]) );
  XOR2X1 U42 ( .A(carry[5]), .B(A[5]), .Y(SUM[5]) );
  AND2X1 U43 ( .A(A[3]), .B(A[4]), .Y(carry[5]) );
  XOR2X1 U44 ( .A(A[3]), .B(A[4]), .Y(SUM[4]) );
endmodule


module Processing_logic_DW01_inc_0 ( A, SUM );
  input [12:0] A;
  output [12:0] SUM;

  wire   [12:2] carry;

  HAX1 U1_1_11 ( .A(A[11]), .B(carry[11]), .YC(carry[12]), .YS(SUM[11]) );
  HAX1 U1_1_10 ( .A(A[10]), .B(carry[10]), .YC(carry[11]), .YS(SUM[10]) );
  HAX1 U1_1_9 ( .A(A[9]), .B(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  HAX1 U1_1_8 ( .A(A[8]), .B(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  HAX1 U1_1_7 ( .A(A[7]), .B(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[12]), .B(A[12]), .Y(SUM[12]) );
endmodule


module Processing_logic_DW01_inc_1 ( A, SUM );
  input [25:0] A;
  output [25:0] SUM;

  wire   [25:2] carry;

  HAX1 U1_1_24 ( .A(A[24]), .B(carry[24]), .YC(carry[25]), .YS(SUM[24]) );
  HAX1 U1_1_23 ( .A(A[23]), .B(carry[23]), .YC(carry[24]), .YS(SUM[23]) );
  HAX1 U1_1_22 ( .A(A[22]), .B(carry[22]), .YC(carry[23]), .YS(SUM[22]) );
  HAX1 U1_1_21 ( .A(A[21]), .B(carry[21]), .YC(carry[22]), .YS(SUM[21]) );
  HAX1 U1_1_20 ( .A(A[20]), .B(carry[20]), .YC(carry[21]), .YS(SUM[20]) );
  HAX1 U1_1_19 ( .A(A[19]), .B(carry[19]), .YC(carry[20]), .YS(SUM[19]) );
  HAX1 U1_1_18 ( .A(A[18]), .B(carry[18]), .YC(carry[19]), .YS(SUM[18]) );
  HAX1 U1_1_17 ( .A(A[17]), .B(carry[17]), .YC(carry[18]), .YS(SUM[17]) );
  HAX1 U1_1_16 ( .A(A[16]), .B(carry[16]), .YC(carry[17]), .YS(SUM[16]) );
  HAX1 U1_1_15 ( .A(A[15]), .B(carry[15]), .YC(carry[16]), .YS(SUM[15]) );
  HAX1 U1_1_14 ( .A(A[14]), .B(carry[14]), .YC(carry[15]), .YS(SUM[14]) );
  HAX1 U1_1_13 ( .A(A[13]), .B(carry[13]), .YC(carry[14]), .YS(SUM[13]) );
  HAX1 U1_1_12 ( .A(A[12]), .B(carry[12]), .YC(carry[13]), .YS(SUM[12]) );
  HAX1 U1_1_11 ( .A(A[11]), .B(carry[11]), .YC(carry[12]), .YS(SUM[11]) );
  HAX1 U1_1_10 ( .A(A[10]), .B(carry[10]), .YC(carry[11]), .YS(SUM[10]) );
  HAX1 U1_1_9 ( .A(A[9]), .B(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  HAX1 U1_1_8 ( .A(A[8]), .B(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  HAX1 U1_1_7 ( .A(A[7]), .B(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[25]), .B(A[25]), .Y(SUM[25]) );
endmodule


module Processing_logic_DW01_inc_2 ( A, SUM );
  input [11:0] A;
  output [11:0] SUM;

  wire   [11:2] carry;

  HAX1 U1_1_10 ( .A(A[10]), .B(carry[10]), .YC(carry[11]), .YS(SUM[10]) );
  HAX1 U1_1_9 ( .A(A[9]), .B(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  HAX1 U1_1_8 ( .A(A[8]), .B(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  HAX1 U1_1_7 ( .A(A[7]), .B(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX1 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[11]), .B(A[11]), .Y(SUM[11]) );
endmodule


module Processing_logic ( DATA_get, CMD_get, RETURN_put, RETURN_address, 
        RETURN_data, cs_bar, ras_bar, cas_bar, we_bar, BA, A, DM, DQS_out, 
        DQ_out, ts_con, modify_setting, clk, ck, reset, ready, CMD_empty, 
        CMD_data_out, DATA_data_out, RETURN_full, DQS_in, DQ_in );
  output [25:0] RETURN_address;
  output [15:0] RETURN_data;
  output [2:0] BA;
  output [12:0] A;
  output [1:0] DM;
  output [1:0] DQS_out;
  output [15:0] DQ_out;
  input [33:0] CMD_data_out;
  input [15:0] DATA_data_out;
  input [1:0] DQS_in;
  input [15:0] DQ_in;
  input clk, ck, reset, ready, CMD_empty, RETURN_full;
  output DATA_get, CMD_get, RETURN_put, cs_bar, ras_bar, cas_bar, we_bar,
         ts_con, modify_setting;
  wire   BLOCK_cmd, DM_flag, listen, ATOMIC_cmd, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n275, n276,
         n284, n350, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n648, n759, n760, n762,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n834, n835, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n890, n1064, n1087,
         n1088, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1120, n1144, n1146, n1147, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n485,
         n486, n487, n488, n490, n491, n492, n493, n495, n496, n497, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n510, n512, n514,
         n515, n516, n517, n518, n519, n520, n521, n523, n525, n526, n527,
         n528, n529, n530, n531, n533, n535, n536, n537, n538, n539, n540,
         n541, n543, n545, n546, n547, n548, n549, n550, n551, n553, n555,
         n556, n557, n558, n559, n560, n561, n563, n565, n566, n567, n568,
         n569, n570, n571, n573, n575, n576, n577, n578, n579, n580, n581,
         n583, n585, n586, n613, n614, n615, n616, n617, n619, n621, n622,
         n623, n624, n625, n626, n627, n641, n643, n644, n645, n646, n647,
         n649, n650, n652, n654, n655, n656, n657, n658, n659, n660, n662,
         n664, n665, n666, n667, n668, n669, n670, n672, n674, n675, n676,
         n677, n678, n679, n680, n682, n684, n688, n689, n690, n691, n692,
         n694, n695, n696, n697, n699, n700, n701, n703, n704, n705, n707,
         n709, n712, n713, n714, n717, n718, n719, n721, n726, n727, n729,
         n731, n733, n735, n737, n739, n741, n743, n745, n747, n749, n751,
         n753, n755, n757, n765, n767, n769, n771, n773, n775, n803, n805,
         n807, n809, n811, n812, n813, n816, n817, n818, n819, n821, n822,
         n824, n825, n826, n827, n829, n830, n831, n832, n833, n836, n837,
         n838, n839, n840, n844, n845, n846, n847, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n863, n864,
         n865, n866, n868, n882, n883, n884, n885, n886, n888, n889, n891,
         n892, n893, n894, n895, n896, n897, n901, n903, n904, n905, n906,
         n909, n912, n914, n915, n918, n919, n920, n921, n922, n923, n924,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n945, n946, n947, n948,
         n949, n951, n952, n953, n954, n956, n958, n960, n961, n962, n965,
         n966, n969, n970, n971, n972, n973, n974, n975, n976, n978, n980,
         n982, n984, n986, n988, n989, n991, n994, n995, n996, n997, n999,
         n1000, n1001, n1002, n1004, n1005, n1007, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1022, n1023, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1034, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1052, n1055, n1056,
         n1057, n1059, n1060, n1061, n1062, n1065, n1066, n1068, n1069, n1071,
         n1073, n1076, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1118, n1119, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1145, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1168, n1169, n1170, n1171, n1173, n1174, n1175, n1176, n1177, n1179,
         n1181, n1182, n1184, n1185, n1186, n1187, n1188, n1190, n1191, n1192,
         n1193, n1195, n1196, n1197, n1198, n1201, n1202, n1203, n1204, n1206,
         n1208, n1210, n1211, n1212, n1213, n1214, n1215, n1217, n1218, n1219,
         n1220, n1223, n1224, n1225, n1227, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1253, n1254, n1256, n1257,
         n1258, n1259, n1260, n1263, n1264, n1265, n1266, n1268, n1270, n1271,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1373, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n277, n278, n279,
         n280, n281, n282, n283, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n489, n494, n498, n499, n509, n511, n513, n522,
         n524, n532, n534, n542, n544, n552, n554, n562, n564, n572, n574,
         n582, n584, n618, n620, n640, n642, n651, n653, n661, n663, n671,
         n673, n681, n683, n685, n686, n687, n693, n698, n702, n706, n708,
         n710, n711, n715, n716, n720, n722, n723, n724, n725, n728, n730,
         n732, n734, n736, n738, n740, n742, n744, n746, n748, n750, n752,
         n754, n756, n758, n761, n763, n764, n766, n768, n770, n772, n774,
         n776, n804, n806, n808, n810, n814, n815, n820, n823, n828, n841,
         n842, n843, n848, n862, n867, n887, n898, n899, n900, n902, n907,
         n908, n910, n911, n913, n916, n917, n925, n944, n950, n955, n957,
         n959, n963, n964, n967, n968, n977, n979, n981, n983, n985, n987,
         n990, n992, n993, n998, n1003, n1006, n1008, n1009, n1021, n1024,
         n1033, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1051, n1053,
         n1054, n1058, n1063, n1067, n1070, n1072, n1074, n1075, n1077, n1078,
         n1089, n1156, n1167, n1172, n1178, n1180, n1183, n1189, n1194, n1199,
         n1200, n1205, n1207, n1209, n1216, n1221, n1222, n1226, n1228, n1239,
         n1251, n1252, n1255, n1261, n1262, n1267, n1269, n1272, n1290, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1374, n1375, n1446, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554;
  wire   [25:3] CMD_addr;
  wire   [12:0] refresh_counter;
  wire   [2:0] state;
  wire   [11:0] counter;
  wire   [1:0] CMD_sz;
  wire   [15:0] ATOMIC_data;
  wire   [2:0] CMD_op;
  wire   [2:0] read_pointer;
  assign cs_bar = 1'b0;

  DFFPOSX1 cas_bar_reg ( .D(n444), .CLK(clk), .Q(cas_bar) );
  DFFPOSX1 ras_bar_reg ( .D(n466), .CLK(clk), .Q(ras_bar) );
  DFFPOSX1 counter_reg_0_ ( .D(n1464), .CLK(clk), .Q(counter[0]) );
  DFFPOSX1 refresh_counter_reg_11_ ( .D(n1359), .CLK(clk), .Q(
        refresh_counter[11]) );
  DFFPOSX1 refresh_counter_reg_12_ ( .D(n1463), .CLK(clk), .Q(
        refresh_counter[12]) );
  DFFPOSX1 CMD_get_reg ( .D(n1444), .CLK(clk), .Q(CMD_get) );
  DFFPOSX1 state_reg_1_ ( .D(n1461), .CLK(clk), .Q(state[1]) );
  DFFPOSX1 ATOMIC_cmd_reg ( .D(n1442), .CLK(clk), .Q(ATOMIC_cmd) );
  DFFPOSX1 BLOCK_cmd_reg ( .D(n1443), .CLK(clk), .Q(BLOCK_cmd) );
  DFFPOSX1 state_reg_2_ ( .D(n1460), .CLK(clk), .Q(state[2]) );
  DFFPOSX1 state_reg_0_ ( .D(n63), .CLK(clk), .Q(state[0]) );
  DFFPOSX1 counter_reg_11_ ( .D(n1445), .CLK(clk), .Q(counter[11]) );
  DFFPOSX1 counter_reg_10_ ( .D(n1447), .CLK(clk), .Q(counter[10]) );
  DFFPOSX1 counter_reg_9_ ( .D(n1448), .CLK(clk), .Q(counter[9]) );
  DFFPOSX1 counter_reg_8_ ( .D(n1449), .CLK(clk), .Q(counter[8]) );
  DFFPOSX1 counter_reg_7_ ( .D(n1450), .CLK(clk), .Q(counter[7]) );
  DFFPOSX1 counter_reg_6_ ( .D(n1451), .CLK(clk), .Q(counter[6]) );
  DFFPOSX1 counter_reg_5_ ( .D(n1452), .CLK(clk), .Q(counter[5]) );
  DFFPOSX1 counter_reg_4_ ( .D(n1453), .CLK(clk), .Q(counter[4]) );
  DFFPOSX1 counter_reg_3_ ( .D(n1454), .CLK(clk), .Q(counter[3]) );
  DFFPOSX1 counter_reg_2_ ( .D(n1455), .CLK(clk), .Q(counter[2]) );
  DFFPOSX1 counter_reg_1_ ( .D(n1456), .CLK(clk), .Q(counter[1]) );
  DFFPOSX1 refresh_counter_reg_0_ ( .D(n1251), .CLK(clk), .Q(
        refresh_counter[0]) );
  DFFPOSX1 refresh_counter_reg_1_ ( .D(n1252), .CLK(clk), .Q(
        refresh_counter[1]) );
  DFFPOSX1 refresh_counter_reg_2_ ( .D(n1255), .CLK(clk), .Q(
        refresh_counter[2]) );
  DFFPOSX1 refresh_counter_reg_3_ ( .D(n1261), .CLK(clk), .Q(
        refresh_counter[3]) );
  DFFPOSX1 refresh_counter_reg_4_ ( .D(n1262), .CLK(clk), .Q(
        refresh_counter[4]) );
  DFFPOSX1 refresh_counter_reg_5_ ( .D(n1267), .CLK(clk), .Q(
        refresh_counter[5]) );
  DFFPOSX1 refresh_counter_reg_6_ ( .D(n1269), .CLK(clk), .Q(
        refresh_counter[6]) );
  DFFPOSX1 refresh_counter_reg_7_ ( .D(n1272), .CLK(clk), .Q(
        refresh_counter[7]) );
  DFFPOSX1 refresh_counter_reg_8_ ( .D(n1290), .CLK(clk), .Q(
        refresh_counter[8]) );
  DFFPOSX1 refresh_counter_reg_9_ ( .D(n1357), .CLK(clk), .Q(
        refresh_counter[9]) );
  DFFPOSX1 refresh_counter_reg_10_ ( .D(n1358), .CLK(clk), .Q(
        refresh_counter[10]) );
  DFFPOSX1 CMD_op_reg_0_ ( .D(n1459), .CLK(clk), .Q(CMD_op[0]) );
  DFFPOSX1 CMD_op_reg_1_ ( .D(n1458), .CLK(clk), .Q(CMD_op[1]) );
  DFFPOSX1 CMD_op_reg_2_ ( .D(n1457), .CLK(clk), .Q(CMD_op[2]) );
  DFFPOSX1 modify_setting_reg ( .D(n449), .CLK(clk), .Q(modify_setting) );
  DFFPOSX1 ts_con_reg ( .D(n65), .CLK(clk), .Q(ts_con) );
  DFFPOSX1 DQS_out_reg_0_ ( .D(n1409), .CLK(clk), .Q(DQS_out[0]) );
  DFFPOSX1 DQS_out_reg_1_ ( .D(n1410), .CLK(clk), .Q(DQS_out[1]) );
  DFFPOSX1 we_bar_reg ( .D(n1222), .CLK(clk), .Q(we_bar) );
  DFFPOSX1 CMD_sz_reg_0_ ( .D(n1414), .CLK(clk), .Q(CMD_sz[0]) );
  DFFPOSX1 CMD_sz_reg_1_ ( .D(n1415), .CLK(clk), .Q(CMD_sz[1]) );
  DFFPOSX1 listen_reg ( .D(n438), .CLK(clk), .Q(listen) );
  DFFPOSX1 DATA_get_reg ( .D(n66), .CLK(clk), .Q(DATA_get) );
  DFFPOSX1 CMD_addr_reg_25_ ( .D(n683), .CLK(clk), .Q(CMD_addr[25]) );
  DFFPOSX1 RETURN_address_reg_25_ ( .D(n1355), .CLK(clk), .Q(
        RETURN_address[25]) );
  DFFPOSX1 CMD_addr_reg_24_ ( .D(n471), .CLK(clk), .Q(CMD_addr[24]) );
  DFFPOSX1 RETURN_address_reg_24_ ( .D(n1354), .CLK(clk), .Q(
        RETURN_address[24]) );
  DFFPOSX1 CMD_addr_reg_0_ ( .D(n446), .CLK(clk), .Q(n759) );
  DFFPOSX1 RETURN_address_reg_0_ ( .D(n1353), .CLK(clk), .Q(RETURN_address[0])
         );
  DFFPOSX1 CMD_addr_reg_1_ ( .D(n309), .CLK(clk), .Q(n760) );
  DFFPOSX1 RETURN_address_reg_1_ ( .D(n1352), .CLK(clk), .Q(RETURN_address[1])
         );
  DFFPOSX1 CMD_addr_reg_2_ ( .D(n318), .CLK(clk), .Q(n762) );
  DFFPOSX1 RETURN_address_reg_2_ ( .D(n1351), .CLK(clk), .Q(RETURN_address[2])
         );
  DFFPOSX1 DM_flag_reg ( .D(n1392), .CLK(clk), .Q(DM_flag) );
  DFFPOSX1 CMD_addr_reg_3_ ( .D(n468), .CLK(clk), .Q(CMD_addr[3]) );
  DFFPOSX1 RETURN_address_reg_3_ ( .D(n1350), .CLK(clk), .Q(RETURN_address[3])
         );
  DFFPOSX1 CMD_addr_reg_4_ ( .D(n327), .CLK(clk), .Q(CMD_addr[4]) );
  DFFPOSX1 RETURN_address_reg_4_ ( .D(n1349), .CLK(clk), .Q(RETURN_address[4])
         );
  DFFPOSX1 CMD_addr_reg_5_ ( .D(n336), .CLK(clk), .Q(CMD_addr[5]) );
  DFFPOSX1 RETURN_address_reg_5_ ( .D(n1348), .CLK(clk), .Q(RETURN_address[5])
         );
  DFFPOSX1 CMD_addr_reg_6_ ( .D(n345), .CLK(clk), .Q(CMD_addr[6]) );
  DFFPOSX1 RETURN_address_reg_6_ ( .D(n1347), .CLK(clk), .Q(RETURN_address[6])
         );
  DFFPOSX1 CMD_addr_reg_7_ ( .D(n357), .CLK(clk), .Q(CMD_addr[7]) );
  DFFPOSX1 RETURN_address_reg_7_ ( .D(n1346), .CLK(clk), .Q(RETURN_address[7])
         );
  DFFPOSX1 CMD_addr_reg_8_ ( .D(n369), .CLK(clk), .Q(CMD_addr[8]) );
  DFFPOSX1 RETURN_address_reg_8_ ( .D(n1345), .CLK(clk), .Q(RETURN_address[8])
         );
  DFFPOSX1 CMD_addr_reg_9_ ( .D(n385), .CLK(clk), .Q(CMD_addr[9]) );
  DFFPOSX1 RETURN_address_reg_9_ ( .D(n1344), .CLK(clk), .Q(RETURN_address[9])
         );
  DFFPOSX1 CMD_addr_reg_10_ ( .D(n400), .CLK(clk), .Q(CMD_addr[10]) );
  DFFPOSX1 RETURN_address_reg_10_ ( .D(n1343), .CLK(clk), .Q(
        RETURN_address[10]) );
  DFFPOSX1 A_reg_0_ ( .D(n67), .CLK(clk), .Q(A[0]) );
  DFFPOSX1 CMD_addr_reg_11_ ( .D(n421), .CLK(clk), .Q(CMD_addr[11]) );
  DFFPOSX1 RETURN_address_reg_11_ ( .D(n1342), .CLK(clk), .Q(
        RETURN_address[11]) );
  DFFPOSX1 A_reg_1_ ( .D(n68), .CLK(clk), .Q(A[1]) );
  DFFPOSX1 CMD_addr_reg_12_ ( .D(n312), .CLK(clk), .Q(CMD_addr[12]) );
  DFFPOSX1 RETURN_address_reg_12_ ( .D(n1341), .CLK(clk), .Q(
        RETURN_address[12]) );
  DFFPOSX1 A_reg_2_ ( .D(n69), .CLK(clk), .Q(A[2]) );
  DFFPOSX1 CMD_addr_reg_13_ ( .D(n321), .CLK(clk), .Q(CMD_addr[13]) );
  DFFPOSX1 RETURN_address_reg_13_ ( .D(n1340), .CLK(clk), .Q(
        RETURN_address[13]) );
  DFFPOSX1 A_reg_3_ ( .D(n70), .CLK(clk), .Q(A[3]) );
  DFFPOSX1 CMD_addr_reg_14_ ( .D(n330), .CLK(clk), .Q(CMD_addr[14]) );
  DFFPOSX1 RETURN_address_reg_14_ ( .D(n1339), .CLK(clk), .Q(
        RETURN_address[14]) );
  DFFPOSX1 A_reg_4_ ( .D(n71), .CLK(clk), .Q(A[4]) );
  DFFPOSX1 CMD_addr_reg_15_ ( .D(n339), .CLK(clk), .Q(CMD_addr[15]) );
  DFFPOSX1 RETURN_address_reg_15_ ( .D(n1338), .CLK(clk), .Q(
        RETURN_address[15]) );
  DFFPOSX1 A_reg_5_ ( .D(n72), .CLK(clk), .Q(A[5]) );
  DFFPOSX1 CMD_addr_reg_16_ ( .D(n348), .CLK(clk), .Q(CMD_addr[16]) );
  DFFPOSX1 RETURN_address_reg_16_ ( .D(n1337), .CLK(clk), .Q(
        RETURN_address[16]) );
  DFFPOSX1 A_reg_6_ ( .D(n73), .CLK(clk), .Q(A[6]) );
  DFFPOSX1 CMD_addr_reg_17_ ( .D(n360), .CLK(clk), .Q(CMD_addr[17]) );
  DFFPOSX1 RETURN_address_reg_17_ ( .D(n1336), .CLK(clk), .Q(
        RETURN_address[17]) );
  DFFPOSX1 A_reg_7_ ( .D(n74), .CLK(clk), .Q(A[7]) );
  DFFPOSX1 CMD_addr_reg_18_ ( .D(n372), .CLK(clk), .Q(CMD_addr[18]) );
  DFFPOSX1 RETURN_address_reg_18_ ( .D(n1335), .CLK(clk), .Q(
        RETURN_address[18]) );
  DFFPOSX1 A_reg_8_ ( .D(n75), .CLK(clk), .Q(A[8]) );
  DFFPOSX1 CMD_addr_reg_19_ ( .D(n388), .CLK(clk), .Q(CMD_addr[19]) );
  DFFPOSX1 RETURN_address_reg_19_ ( .D(n1334), .CLK(clk), .Q(
        RETURN_address[19]) );
  DFFPOSX1 A_reg_9_ ( .D(n76), .CLK(clk), .Q(A[9]) );
  DFFPOSX1 CMD_addr_reg_20_ ( .D(n403), .CLK(clk), .Q(CMD_addr[20]) );
  DFFPOSX1 RETURN_address_reg_20_ ( .D(n1333), .CLK(clk), .Q(
        RETURN_address[20]) );
  DFFPOSX1 A_reg_10_ ( .D(n1221), .CLK(clk), .Q(A[10]) );
  DFFPOSX1 CMD_addr_reg_21_ ( .D(n424), .CLK(clk), .Q(CMD_addr[21]) );
  DFFPOSX1 RETURN_address_reg_21_ ( .D(n1332), .CLK(clk), .Q(
        RETURN_address[21]) );
  DFFPOSX1 A_reg_11_ ( .D(n1396), .CLK(clk), .Q(A[11]) );
  DFFPOSX1 CMD_addr_reg_22_ ( .D(n441), .CLK(clk), .Q(CMD_addr[22]) );
  DFFPOSX1 RETURN_address_reg_22_ ( .D(n1331), .CLK(clk), .Q(
        RETURN_address[22]) );
  DFFPOSX1 A_reg_12_ ( .D(n1395), .CLK(clk), .Q(A[12]) );
  DFFPOSX1 CMD_addr_reg_23_ ( .D(n687), .CLK(clk), .Q(CMD_addr[23]) );
  DFFPOSX1 RETURN_address_reg_23_ ( .D(n1330), .CLK(clk), .Q(
        RETURN_address[23]) );
  DFFPOSX1 BA_reg_0_ ( .D(n77), .CLK(clk), .Q(BA[0]) );
  DFFPOSX1 BA_reg_1_ ( .D(n1394), .CLK(clk), .Q(BA[1]) );
  DFFPOSX1 BA_reg_2_ ( .D(n1393), .CLK(clk), .Q(BA[2]) );
  DFFPOSX1 read_pointer_reg_0_ ( .D(n1329), .CLK(clk), .Q(read_pointer[0]) );
  DFFPOSX1 read_pointer_reg_1_ ( .D(n1328), .CLK(clk), .Q(read_pointer[1]) );
  DFFPOSX1 read_pointer_reg_2_ ( .D(n1327), .CLK(clk), .Q(read_pointer[2]) );
  DFFPOSX1 ATOMIC_data_reg_0_ ( .D(n2), .CLK(clk), .Q(ATOMIC_data[0]) );
  DFFPOSX1 ATOMIC_data_reg_1_ ( .D(n3), .CLK(clk), .Q(ATOMIC_data[1]) );
  DFFPOSX1 ATOMIC_data_reg_2_ ( .D(n4), .CLK(clk), .Q(ATOMIC_data[2]) );
  DFFPOSX1 ATOMIC_data_reg_3_ ( .D(n5), .CLK(clk), .Q(ATOMIC_data[3]) );
  DFFPOSX1 ATOMIC_data_reg_4_ ( .D(n6), .CLK(clk), .Q(ATOMIC_data[4]) );
  DFFPOSX1 ATOMIC_data_reg_5_ ( .D(n7), .CLK(clk), .Q(ATOMIC_data[5]) );
  DFFPOSX1 ATOMIC_data_reg_6_ ( .D(n8), .CLK(clk), .Q(ATOMIC_data[6]) );
  DFFPOSX1 ATOMIC_data_reg_8_ ( .D(n9), .CLK(clk), .Q(ATOMIC_data[8]) );
  DFFPOSX1 ATOMIC_data_reg_9_ ( .D(n10), .CLK(clk), .Q(ATOMIC_data[9]) );
  DFFPOSX1 ATOMIC_data_reg_10_ ( .D(n11), .CLK(clk), .Q(ATOMIC_data[10]) );
  DFFPOSX1 ATOMIC_data_reg_11_ ( .D(n12), .CLK(clk), .Q(ATOMIC_data[11]) );
  DFFPOSX1 ATOMIC_data_reg_12_ ( .D(n13), .CLK(clk), .Q(ATOMIC_data[12]) );
  DFFPOSX1 ATOMIC_data_reg_13_ ( .D(n14), .CLK(clk), .Q(ATOMIC_data[13]) );
  DFFPOSX1 ATOMIC_data_reg_14_ ( .D(n15), .CLK(clk), .Q(ATOMIC_data[14]) );
  DFFPOSX1 ATOMIC_data_reg_7_ ( .D(n16), .CLK(clk), .Q(ATOMIC_data[7]) );
  DFFPOSX1 ATOMIC_data_reg_15_ ( .D(n17), .CLK(clk), .Q(ATOMIC_data[15]) );
  DFFPOSX1 RETURN_put_reg ( .D(n64), .CLK(clk), .Q(RETURN_put) );
  DFFNEGX1 DM_reg_1_ ( .D(n1510), .CLK(clk), .Q(DM[1]) );
  DFFNEGX1 DM_reg_0_ ( .D(n1510), .CLK(clk), .Q(DM[0]) );
  DFFNEGX1 DQ_out_reg_15_ ( .D(n1391), .CLK(clk), .Q(DQ_out[15]) );
  DFFNEGX1 DQ_out_reg_14_ ( .D(n1390), .CLK(clk), .Q(DQ_out[14]) );
  DFFNEGX1 DQ_out_reg_13_ ( .D(n1389), .CLK(clk), .Q(DQ_out[13]) );
  DFFNEGX1 DQ_out_reg_12_ ( .D(n1388), .CLK(clk), .Q(DQ_out[12]) );
  DFFNEGX1 DQ_out_reg_11_ ( .D(n1387), .CLK(clk), .Q(DQ_out[11]) );
  DFFNEGX1 DQ_out_reg_10_ ( .D(n1386), .CLK(clk), .Q(DQ_out[10]) );
  DFFNEGX1 DQ_out_reg_9_ ( .D(n1385), .CLK(clk), .Q(DQ_out[9]) );
  DFFNEGX1 DQ_out_reg_8_ ( .D(n1384), .CLK(clk), .Q(DQ_out[8]) );
  DFFNEGX1 DQ_out_reg_7_ ( .D(n1383), .CLK(clk), .Q(DQ_out[7]) );
  DFFNEGX1 DQ_out_reg_6_ ( .D(n1382), .CLK(clk), .Q(DQ_out[6]) );
  DFFNEGX1 DQ_out_reg_5_ ( .D(n1381), .CLK(clk), .Q(DQ_out[5]) );
  DFFNEGX1 DQ_out_reg_4_ ( .D(n1380), .CLK(clk), .Q(DQ_out[4]) );
  DFFNEGX1 DQ_out_reg_3_ ( .D(n1379), .CLK(clk), .Q(DQ_out[3]) );
  DFFNEGX1 DQ_out_reg_2_ ( .D(n1378), .CLK(clk), .Q(DQ_out[2]) );
  DFFNEGX1 DQ_out_reg_1_ ( .D(n1377), .CLK(clk), .Q(DQ_out[1]) );
  DFFNEGX1 DQ_out_reg_0_ ( .D(n1376), .CLK(clk), .Q(DQ_out[0]) );
  NAND3X1 U3 ( .A(n202), .B(n237), .C(n256), .Y(n1295) );
  AOI21X1 U5 ( .A(reset), .B(ATOMIC_data[15]), .C(n488), .Y(n487) );
  OAI21X1 U6 ( .A(n1553), .B(n483), .C(n142), .Y(n488) );
  AOI22X1 U8 ( .A(n493), .B(n1070), .C(RETURN_data[15]), .D(n495), .Y(n486) );
  OAI21X1 U9 ( .A(n1553), .B(n1035), .C(n137), .Y(n495) );
  AOI21X1 U10 ( .A(n1496), .B(n1553), .C(n1037), .Y(n497) );
  OAI21X1 U12 ( .A(n459), .B(n1553), .C(n501), .Y(n493) );
  AOI22X1 U13 ( .A(RETURN_data[14]), .B(n502), .C(n503), .D(n1325), .Y(n485)
         );
  NAND3X1 U14 ( .A(n201), .B(n236), .C(n506), .Y(n1296) );
  AOI22X1 U16 ( .A(n1021), .B(RETURN_data[15]), .C(DATA_data_out[7]), .D(n1037), .Y(n508) );
  AOI22X1 U17 ( .A(RETURN_data[8]), .B(n1495), .C(ATOMIC_data[7]), .D(reset), 
        .Y(n507) );
  AOI22X1 U18 ( .A(n510), .B(n1167), .C(RETURN_data[7]), .D(n512), .Y(n505) );
  OAI21X1 U19 ( .A(n1035), .B(n1545), .C(n136), .Y(n512) );
  AOI21X1 U20 ( .A(n1496), .B(n1545), .C(n1037), .Y(n514) );
  OAI21X1 U23 ( .A(n1036), .B(n1545), .C(n501), .Y(n510) );
  AOI22X1 U26 ( .A(RETURN_data[6]), .B(n502), .C(n1317), .D(n503), .Y(n504) );
  NAND3X1 U27 ( .A(n200), .B(n235), .C(n518), .Y(n1297) );
  AOI22X1 U30 ( .A(RETURN_data[6]), .B(n1024), .C(DATA_data_out[14]), .D(n1037), .Y(n520) );
  AOI22X1 U31 ( .A(n1495), .B(RETURN_data[15]), .C(ATOMIC_data[14]), .D(reset), 
        .Y(n519) );
  AOI22X1 U32 ( .A(n521), .B(n1072), .C(RETURN_data[14]), .D(n523), .Y(n517)
         );
  OAI21X1 U33 ( .A(n1035), .B(n1552), .C(n135), .Y(n523) );
  AOI21X1 U34 ( .A(n1496), .B(n1552), .C(n1037), .Y(n525) );
  OAI21X1 U36 ( .A(n1036), .B(n1552), .C(n501), .Y(n521) );
  AOI22X1 U37 ( .A(RETURN_data[13]), .B(n502), .C(n1324), .D(n503), .Y(n516)
         );
  NAND3X1 U38 ( .A(n199), .B(n234), .C(n528), .Y(n1298) );
  AOI22X1 U40 ( .A(RETURN_data[5]), .B(n1024), .C(DATA_data_out[13]), .D(n1037), .Y(n530) );
  AOI22X1 U41 ( .A(n1495), .B(RETURN_data[14]), .C(ATOMIC_data[13]), .D(reset), 
        .Y(n529) );
  AOI22X1 U42 ( .A(n531), .B(n1074), .C(RETURN_data[13]), .D(n533), .Y(n527)
         );
  OAI21X1 U43 ( .A(n1035), .B(n1551), .C(n134), .Y(n533) );
  AOI21X1 U44 ( .A(n1496), .B(n1551), .C(n1037), .Y(n535) );
  OAI21X1 U46 ( .A(n1036), .B(n1551), .C(n501), .Y(n531) );
  AOI22X1 U47 ( .A(RETURN_data[12]), .B(n502), .C(n1323), .D(n503), .Y(n526)
         );
  NAND3X1 U48 ( .A(n198), .B(n233), .C(n538), .Y(n1299) );
  AOI22X1 U50 ( .A(RETURN_data[4]), .B(n1024), .C(DATA_data_out[12]), .D(n1037), .Y(n540) );
  AOI22X1 U51 ( .A(RETURN_data[13]), .B(n1495), .C(ATOMIC_data[12]), .D(reset), 
        .Y(n539) );
  AOI22X1 U52 ( .A(n541), .B(n1075), .C(RETURN_data[12]), .D(n543), .Y(n537)
         );
  OAI21X1 U53 ( .A(n1035), .B(n1550), .C(n133), .Y(n543) );
  AOI21X1 U54 ( .A(n1496), .B(n1550), .C(n1037), .Y(n545) );
  OAI21X1 U56 ( .A(n1036), .B(n1550), .C(n501), .Y(n541) );
  AOI22X1 U57 ( .A(RETURN_data[11]), .B(n502), .C(n1322), .D(n503), .Y(n536)
         );
  NAND3X1 U58 ( .A(n197), .B(n232), .C(n548), .Y(n1300) );
  AOI22X1 U60 ( .A(RETURN_data[3]), .B(n1024), .C(DATA_data_out[11]), .D(n1037), .Y(n550) );
  AOI22X1 U61 ( .A(RETURN_data[12]), .B(n1495), .C(ATOMIC_data[11]), .D(reset), 
        .Y(n549) );
  AOI22X1 U62 ( .A(n551), .B(n1077), .C(RETURN_data[11]), .D(n553), .Y(n547)
         );
  OAI21X1 U63 ( .A(n1035), .B(n1549), .C(n132), .Y(n553) );
  AOI21X1 U64 ( .A(n1496), .B(n1549), .C(n1037), .Y(n555) );
  OAI21X1 U66 ( .A(n1036), .B(n1549), .C(n501), .Y(n551) );
  AOI22X1 U67 ( .A(RETURN_data[10]), .B(n502), .C(n1321), .D(n503), .Y(n546)
         );
  NAND3X1 U68 ( .A(n196), .B(n231), .C(n558), .Y(n1301) );
  AOI22X1 U70 ( .A(RETURN_data[2]), .B(n1024), .C(DATA_data_out[10]), .D(n1037), .Y(n560) );
  AOI22X1 U71 ( .A(RETURN_data[11]), .B(n1495), .C(ATOMIC_data[10]), .D(reset), 
        .Y(n559) );
  AOI22X1 U72 ( .A(n561), .B(n1078), .C(RETURN_data[10]), .D(n563), .Y(n557)
         );
  OAI21X1 U73 ( .A(n1035), .B(n1548), .C(n131), .Y(n563) );
  AOI21X1 U74 ( .A(n1496), .B(n1548), .C(n1037), .Y(n565) );
  OAI21X1 U76 ( .A(n1036), .B(n1548), .C(n501), .Y(n561) );
  AOI22X1 U77 ( .A(RETURN_data[9]), .B(n502), .C(n1320), .D(n503), .Y(n556) );
  NAND3X1 U78 ( .A(n195), .B(n230), .C(n568), .Y(n1302) );
  AOI22X1 U80 ( .A(RETURN_data[1]), .B(n1024), .C(DATA_data_out[9]), .D(n1037), 
        .Y(n570) );
  AOI22X1 U81 ( .A(RETURN_data[10]), .B(n1495), .C(ATOMIC_data[9]), .D(reset), 
        .Y(n569) );
  AOI22X1 U82 ( .A(n571), .B(n1089), .C(RETURN_data[9]), .D(n573), .Y(n567) );
  OAI21X1 U83 ( .A(n1035), .B(n1547), .C(n130), .Y(n573) );
  AOI21X1 U84 ( .A(n1496), .B(n1547), .C(n1037), .Y(n575) );
  OAI21X1 U86 ( .A(n1036), .B(n1547), .C(n501), .Y(n571) );
  AOI22X1 U87 ( .A(RETURN_data[8]), .B(n502), .C(n1319), .D(n503), .Y(n566) );
  NAND3X1 U88 ( .A(n194), .B(n229), .C(n578), .Y(n1303) );
  AOI22X1 U90 ( .A(RETURN_data[0]), .B(n1024), .C(DATA_data_out[8]), .D(n1037), 
        .Y(n580) );
  AOI22X1 U91 ( .A(RETURN_data[9]), .B(n1495), .C(ATOMIC_data[8]), .D(reset), 
        .Y(n579) );
  AOI22X1 U92 ( .A(n581), .B(n1156), .C(RETURN_data[8]), .D(n583), .Y(n577) );
  OAI21X1 U93 ( .A(n1035), .B(n1546), .C(n129), .Y(n583) );
  AOI21X1 U94 ( .A(n1496), .B(n1546), .C(n1037), .Y(n585) );
  OAI21X1 U96 ( .A(n1036), .B(n1546), .C(n501), .Y(n581) );
  AOI22X1 U97 ( .A(RETURN_data[7]), .B(n502), .C(n1318), .D(n503), .Y(n576) );
  NAND3X1 U98 ( .A(n193), .B(n228), .C(n614), .Y(n1304) );
  AOI22X1 U100 ( .A(n1021), .B(RETURN_data[14]), .C(DATA_data_out[6]), .D(
        n1037), .Y(n616) );
  AOI22X1 U101 ( .A(n1495), .B(RETURN_data[7]), .C(ATOMIC_data[6]), .D(reset), 
        .Y(n615) );
  AOI22X1 U102 ( .A(n617), .B(n1172), .C(RETURN_data[6]), .D(n619), .Y(n613)
         );
  OAI21X1 U103 ( .A(n1035), .B(n1544), .C(n128), .Y(n619) );
  AOI21X1 U104 ( .A(n1496), .B(n1544), .C(n1037), .Y(n621) );
  OAI21X1 U106 ( .A(n1036), .B(n1544), .C(n501), .Y(n617) );
  AOI22X1 U107 ( .A(RETURN_data[5]), .B(n502), .C(n1316), .D(n503), .Y(n586)
         );
  NAND3X1 U108 ( .A(n192), .B(n227), .C(n624), .Y(n1305) );
  AOI22X1 U110 ( .A(RETURN_data[13]), .B(n1021), .C(DATA_data_out[5]), .D(
        n1037), .Y(n626) );
  AOI22X1 U111 ( .A(n1495), .B(RETURN_data[6]), .C(ATOMIC_data[5]), .D(reset), 
        .Y(n625) );
  AOI22X1 U112 ( .A(n627), .B(n1178), .C(RETURN_data[5]), .D(n641), .Y(n623)
         );
  OAI21X1 U113 ( .A(n1035), .B(n1543), .C(n127), .Y(n641) );
  AOI21X1 U114 ( .A(n1496), .B(n1543), .C(n1037), .Y(n643) );
  OAI21X1 U116 ( .A(n1036), .B(n1543), .C(n501), .Y(n627) );
  AOI22X1 U117 ( .A(RETURN_data[4]), .B(n502), .C(n1315), .D(n503), .Y(n622)
         );
  NAND3X1 U118 ( .A(n191), .B(n226), .C(n646), .Y(n1306) );
  AOI22X1 U120 ( .A(RETURN_data[12]), .B(n1021), .C(DATA_data_out[4]), .D(
        n1037), .Y(n649) );
  AOI22X1 U121 ( .A(RETURN_data[5]), .B(n1495), .C(ATOMIC_data[4]), .D(reset), 
        .Y(n647) );
  AOI22X1 U122 ( .A(n650), .B(n1180), .C(RETURN_data[4]), .D(n652), .Y(n645)
         );
  OAI21X1 U123 ( .A(n1035), .B(n1542), .C(n126), .Y(n652) );
  AOI21X1 U124 ( .A(n1496), .B(n1542), .C(n1037), .Y(n654) );
  OAI21X1 U126 ( .A(n1036), .B(n1542), .C(n501), .Y(n650) );
  AOI22X1 U127 ( .A(RETURN_data[3]), .B(n502), .C(n1314), .D(n503), .Y(n644)
         );
  NAND3X1 U128 ( .A(n190), .B(n225), .C(n657), .Y(n1307) );
  AOI22X1 U130 ( .A(RETURN_data[11]), .B(n1021), .C(DATA_data_out[3]), .D(
        n1037), .Y(n659) );
  AOI22X1 U131 ( .A(RETURN_data[4]), .B(n1495), .C(ATOMIC_data[3]), .D(reset), 
        .Y(n658) );
  AOI22X1 U132 ( .A(n660), .B(n1183), .C(RETURN_data[3]), .D(n662), .Y(n656)
         );
  OAI21X1 U133 ( .A(n1035), .B(n1541), .C(n125), .Y(n662) );
  AOI21X1 U134 ( .A(n1496), .B(n1541), .C(n1037), .Y(n664) );
  OAI21X1 U136 ( .A(n1036), .B(n1541), .C(n501), .Y(n660) );
  AOI22X1 U137 ( .A(RETURN_data[2]), .B(n502), .C(n1313), .D(n503), .Y(n655)
         );
  NAND3X1 U138 ( .A(n189), .B(n224), .C(n667), .Y(n1308) );
  AOI22X1 U140 ( .A(RETURN_data[10]), .B(n1021), .C(DATA_data_out[2]), .D(
        n1037), .Y(n669) );
  AOI22X1 U141 ( .A(RETURN_data[3]), .B(n1495), .C(ATOMIC_data[2]), .D(reset), 
        .Y(n668) );
  AOI22X1 U142 ( .A(n670), .B(n1189), .C(RETURN_data[2]), .D(n672), .Y(n666)
         );
  OAI21X1 U143 ( .A(n1035), .B(n1540), .C(n124), .Y(n672) );
  AOI21X1 U144 ( .A(n1496), .B(n1540), .C(n1037), .Y(n674) );
  OAI21X1 U146 ( .A(n1036), .B(n1540), .C(n501), .Y(n670) );
  AOI22X1 U147 ( .A(RETURN_data[1]), .B(n502), .C(n1312), .D(n503), .Y(n665)
         );
  NAND3X1 U148 ( .A(n188), .B(n223), .C(n677), .Y(n1309) );
  AOI22X1 U150 ( .A(RETURN_data[9]), .B(n1021), .C(DATA_data_out[1]), .D(n1037), .Y(n679) );
  AOI22X1 U151 ( .A(RETURN_data[2]), .B(n1495), .C(ATOMIC_data[1]), .D(reset), 
        .Y(n678) );
  AOI22X1 U152 ( .A(n680), .B(n1194), .C(RETURN_data[1]), .D(n682), .Y(n676)
         );
  OAI21X1 U153 ( .A(n1035), .B(n1539), .C(n123), .Y(n682) );
  AOI21X1 U154 ( .A(n1496), .B(n1539), .C(n1037), .Y(n684) );
  OAI21X1 U156 ( .A(n1036), .B(n1539), .C(n501), .Y(n680) );
  NAND3X1 U157 ( .A(n1498), .B(n1063), .C(n1497), .Y(n515) );
  AOI22X1 U158 ( .A(RETURN_data[0]), .B(n502), .C(n1311), .D(n503), .Y(n675)
         );
  NAND3X1 U160 ( .A(n187), .B(n222), .C(n255), .Y(n1326) );
  AOI21X1 U161 ( .A(ATOMIC_data[0]), .B(reset), .C(n692), .Y(n691) );
  OAI21X1 U162 ( .A(n483), .B(n1538), .C(n141), .Y(n692) );
  NAND3X1 U165 ( .A(CMD_op[1]), .B(CMD_op[2]), .C(n696), .Y(n695) );
  AOI22X1 U167 ( .A(n697), .B(n1199), .C(RETURN_data[0]), .D(n699), .Y(n690)
         );
  OAI21X1 U168 ( .A(n1035), .B(n1538), .C(n122), .Y(n699) );
  AOI21X1 U169 ( .A(n1496), .B(n1538), .C(n1037), .Y(n700) );
  NAND3X1 U171 ( .A(CMD_op[1]), .B(n1497), .C(n701), .Y(n490) );
  NAND3X1 U174 ( .A(n1499), .B(n1063), .C(CMD_op[1]), .Y(n496) );
  OAI21X1 U176 ( .A(n459), .B(n1538), .C(n501), .Y(n697) );
  NAND3X1 U178 ( .A(CMD_op[2]), .B(n1497), .C(n704), .Y(n500) );
  AOI22X1 U180 ( .A(n1310), .B(n503), .C(RETURN_data[8]), .D(n1021), .Y(n689)
         );
  NOR3X1 U182 ( .A(n1499), .B(reset), .C(n1497), .Y(n688) );
  NOR3X1 U184 ( .A(CMD_op[2]), .B(reset), .C(CMD_op[1]), .Y(n703) );
  OAI21X1 U185 ( .A(n451), .B(n1534), .C(n452), .Y(n1327) );
  NAND3X1 U186 ( .A(n1372), .B(n1534), .C(read_pointer[1]), .Y(n707) );
  AOI21X1 U189 ( .A(n714), .B(n1533), .C(n712), .Y(n705) );
  OAI21X1 U191 ( .A(read_pointer[1]), .B(n477), .C(n419), .Y(n1328) );
  OAI21X1 U193 ( .A(read_pointer[0]), .B(n716), .C(n1374), .Y(n712) );
  NAND3X1 U194 ( .A(n714), .B(n1374), .C(read_pointer[0]), .Y(n709) );
  OAI21X1 U195 ( .A(n1374), .B(n1532), .C(n121), .Y(n1329) );
  NAND3X1 U196 ( .A(n1374), .B(n1532), .C(n714), .Y(n717) );
  NAND3X1 U200 ( .A(n207), .B(n1063), .C(n1476), .Y(n718) );
  NAND3X1 U203 ( .A(n1059), .B(n1026), .C(n726), .Y(n721) );
  OAI21X1 U205 ( .A(reset), .B(n1531), .C(n464), .Y(n1330) );
  OAI21X1 U208 ( .A(reset), .B(n1530), .C(n671), .Y(n1331) );
  OAI21X1 U210 ( .A(reset), .B(n1529), .C(n663), .Y(n1332) );
  OAI21X1 U212 ( .A(reset), .B(n1528), .C(n661), .Y(n1333) );
  OAI21X1 U215 ( .A(reset), .B(n1527), .C(n653), .Y(n1334) );
  OAI21X1 U218 ( .A(reset), .B(n1526), .C(n651), .Y(n1335) );
  OAI21X1 U221 ( .A(reset), .B(n1525), .C(n642), .Y(n1336) );
  OAI21X1 U224 ( .A(reset), .B(n1524), .C(n640), .Y(n1337) );
  OAI21X1 U227 ( .A(reset), .B(n1523), .C(n620), .Y(n1338) );
  OAI21X1 U230 ( .A(reset), .B(n1522), .C(n618), .Y(n1339) );
  OAI21X1 U233 ( .A(reset), .B(n1521), .C(n584), .Y(n1340) );
  OAI21X1 U236 ( .A(reset), .B(n1520), .C(n582), .Y(n1341) );
  OAI21X1 U239 ( .A(reset), .B(n1519), .C(n574), .Y(n1342) );
  OAI21X1 U242 ( .A(reset), .B(n1518), .C(n572), .Y(n1343) );
  OAI21X1 U245 ( .A(reset), .B(n1517), .C(n564), .Y(n1344) );
  OAI21X1 U248 ( .A(reset), .B(n1516), .C(n562), .Y(n1345) );
  OAI21X1 U251 ( .A(reset), .B(n1515), .C(n554), .Y(n1346) );
  OAI21X1 U254 ( .A(reset), .B(n1514), .C(n552), .Y(n1347) );
  OAI21X1 U257 ( .A(reset), .B(n1513), .C(n544), .Y(n1348) );
  OAI21X1 U260 ( .A(reset), .B(n1512), .C(n542), .Y(n1349) );
  OAI21X1 U263 ( .A(reset), .B(n1511), .C(n534), .Y(n1350) );
  OAI21X1 U266 ( .A(reset), .B(n1509), .C(n532), .Y(n1351) );
  OAI21X1 U268 ( .A(reset), .B(n1508), .C(n524), .Y(n1352) );
  OAI21X1 U270 ( .A(reset), .B(n1507), .C(n522), .Y(n1353) );
  OAI21X1 U273 ( .A(reset), .B(n1506), .C(n513), .Y(n1354) );
  OAI21X1 U275 ( .A(reset), .B(n1505), .C(n511), .Y(n1355) );
  AOI22X1 U279 ( .A(n1228), .B(CMD_addr[23]), .C(n288), .D(n817), .Y(n812) );
  AOI22X1 U282 ( .A(n822), .B(n213), .C(A[10]), .D(n289), .Y(n819) );
  NAND3X1 U283 ( .A(n1478), .B(n824), .C(n254), .Y(n821) );
  AOI21X1 U284 ( .A(n304), .B(CMD_addr[20]), .C(n827), .Y(n825) );
  OAI21X1 U285 ( .A(n831), .B(n461), .C(n396), .Y(n827) );
  NAND3X1 U290 ( .A(n291), .B(n241), .C(n249), .Y(n836) );
  AOI22X1 U291 ( .A(n219), .B(n1360), .C(n1361), .D(n995), .Y(n839) );
  AOI21X1 U293 ( .A(n414), .B(n379), .C(n481), .Y(n840) );
  AOI22X1 U296 ( .A(n102), .B(n847), .C(refresh_counter[0]), .D(n860), .Y(n846) );
  AOI22X1 U298 ( .A(n103), .B(n847), .C(refresh_counter[1]), .D(n860), .Y(n849) );
  AOI22X1 U300 ( .A(n104), .B(n847), .C(refresh_counter[2]), .D(n860), .Y(n850) );
  AOI22X1 U302 ( .A(n105), .B(n847), .C(refresh_counter[3]), .D(n860), .Y(n851) );
  AOI22X1 U304 ( .A(n106), .B(n847), .C(refresh_counter[4]), .D(n860), .Y(n852) );
  AOI22X1 U306 ( .A(n107), .B(n847), .C(refresh_counter[5]), .D(n860), .Y(n853) );
  AOI22X1 U308 ( .A(n108), .B(n847), .C(refresh_counter[6]), .D(n860), .Y(n854) );
  AOI22X1 U310 ( .A(n109), .B(n847), .C(refresh_counter[7]), .D(n860), .Y(n855) );
  AOI22X1 U312 ( .A(n110), .B(n847), .C(refresh_counter[8]), .D(n860), .Y(n856) );
  AOI22X1 U314 ( .A(n111), .B(n847), .C(refresh_counter[9]), .D(n860), .Y(n857) );
  AOI22X1 U316 ( .A(n112), .B(n847), .C(refresh_counter[10]), .D(n860), .Y(
        n858) );
  AOI22X1 U318 ( .A(n113), .B(n847), .C(refresh_counter[11]), .D(n860), .Y(
        n859) );
  OAI21X1 U321 ( .A(n1500), .B(n863), .C(ready), .Y(n861) );
  OAI21X1 U323 ( .A(n865), .B(n480), .C(n1360), .Y(n864) );
  OAI21X1 U325 ( .A(n1510), .B(n292), .C(n120), .Y(n1392) );
  NAND3X1 U326 ( .A(n292), .B(n1063), .C(n253), .Y(n868) );
  NAND3X1 U327 ( .A(n482), .B(n725), .C(n248), .Y(n882) );
  AOI22X1 U328 ( .A(n221), .B(n1510), .C(BLOCK_cmd), .D(n1369), .Y(n885) );
  NOR3X1 U331 ( .A(n894), .B(reset), .C(n298), .Y(n893) );
  NOR3X1 U332 ( .A(n264), .B(n759), .C(n265), .Y(n894) );
  AOI22X1 U333 ( .A(n1366), .B(n995), .C(n1365), .D(n1027), .Y(n897) );
  NAND3X1 U338 ( .A(n1027), .B(n901), .C(n1369), .Y(n892) );
  OAI21X1 U340 ( .A(n1), .B(n246), .C(n1510), .Y(n901) );
  NAND3X1 U341 ( .A(n904), .B(n905), .C(n906), .Y(n903) );
  XNOR2X1 U342 ( .A(counter[0]), .B(n759), .Y(n906) );
  XNOR2X1 U344 ( .A(counter[1]), .B(n760), .Y(n904) );
  NAND3X1 U348 ( .A(n995), .B(n909), .C(n1368), .Y(n891) );
  OAI21X1 U350 ( .A(n905), .B(n429), .C(n1510), .Y(n909) );
  NAND3X1 U351 ( .A(n1492), .B(n914), .C(n915), .Y(n912) );
  XNOR2X1 U352 ( .A(counter[0]), .B(n759), .Y(n915) );
  XNOR2X1 U353 ( .A(counter[1]), .B(n760), .Y(n914) );
  OAI21X1 U359 ( .A(n1505), .B(n818), .C(n436), .Y(n1393) );
  OAI21X1 U362 ( .A(n1506), .B(n818), .C(n418), .Y(n1394) );
  OAI21X1 U365 ( .A(n1530), .B(n818), .C(n397), .Y(n1395) );
  OAI21X1 U368 ( .A(n1529), .B(n818), .C(n382), .Y(n1396) );
  AOI22X1 U374 ( .A(n1006), .B(CMD_addr[9]), .C(n1009), .D(CMD_addr[19]), .Y(
        n923) );
  AOI22X1 U376 ( .A(n1006), .B(CMD_addr[8]), .C(n1009), .D(CMD_addr[18]), .Y(
        n929) );
  AOI22X1 U377 ( .A(A[8]), .B(n930), .C(n307), .D(n931), .Y(n928) );
  AOI22X1 U380 ( .A(n1006), .B(CMD_addr[7]), .C(n1009), .D(CMD_addr[17]), .Y(
        n932) );
  AOI22X1 U383 ( .A(n1006), .B(CMD_addr[6]), .C(n1009), .D(CMD_addr[16]), .Y(
        n934) );
  AOI22X1 U386 ( .A(n1006), .B(CMD_addr[5]), .C(n1008), .D(CMD_addr[15]), .Y(
        n936) );
  AOI22X1 U388 ( .A(n220), .B(n307), .C(n1003), .D(CMD_addr[4]), .Y(n939) );
  AOI22X1 U391 ( .A(n1009), .B(CMD_addr[14]), .C(A[4]), .D(n930), .Y(n938) );
  AOI22X1 U393 ( .A(n1003), .B(CMD_addr[3]), .C(n1008), .D(CMD_addr[13]), .Y(
        n943) );
  AOI22X1 U394 ( .A(A[3]), .B(n930), .C(n269), .D(n307), .Y(n942) );
  AOI22X1 U396 ( .A(n1003), .B(n762), .C(n1008), .D(CMD_addr[12]), .Y(n946) );
  AOI22X1 U397 ( .A(A[2]), .B(n930), .C(n269), .D(n307), .Y(n945) );
  AOI22X1 U400 ( .A(n1003), .B(n760), .C(n1008), .D(CMD_addr[11]), .Y(n949) );
  AOI22X1 U401 ( .A(A[1]), .B(n930), .C(n1481), .D(n307), .Y(n948) );
  AOI22X1 U406 ( .A(n1003), .B(n759), .C(n1008), .D(CMD_addr[10]), .Y(n952) );
  NAND3X1 U410 ( .A(n1476), .B(n1063), .C(n302), .Y(n954) );
  AOI21X1 U413 ( .A(n1476), .B(n304), .C(n1239), .Y(n837) );
  NAND3X1 U415 ( .A(n1472), .B(n865), .C(n1360), .Y(n956) );
  OAI21X1 U417 ( .A(n454), .B(n941), .C(n270), .Y(n817) );
  NAND3X1 U418 ( .A(n1164), .B(n960), .C(n961), .Y(n947) );
  OAI21X1 U419 ( .A(n941), .B(n478), .C(n453), .Y(n931) );
  NAND3X1 U420 ( .A(n1059), .B(n1489), .C(n1482), .Y(n951) );
  NAND3X1 U422 ( .A(counter[5]), .B(counter[4]), .C(counter[7]), .Y(n966) );
  NAND3X1 U423 ( .A(n1479), .B(n1487), .C(counter[2]), .Y(n965) );
  AOI21X1 U426 ( .A(n1500), .B(n450), .C(reset), .Y(n1407) );
  NAND3X1 U430 ( .A(n283), .B(n1063), .C(n263), .Y(n972) );
  AOI22X1 U435 ( .A(n1027), .B(n980), .C(n1200), .D(n995), .Y(n978) );
  OAI21X1 U436 ( .A(BLOCK_cmd), .B(n725), .C(n119), .Y(n980) );
  AOI21X1 U437 ( .A(n1012), .B(n984), .C(n1375), .Y(n982) );
  OAI21X1 U439 ( .A(n986), .B(n1501), .C(n118), .Y(n1409) );
  NAND3X1 U440 ( .A(n457), .B(n1501), .C(n986), .Y(n988) );
  OAI21X1 U442 ( .A(n986), .B(n1502), .C(n117), .Y(n1410) );
  NAND3X1 U443 ( .A(n457), .B(n1502), .C(n986), .Y(n991) );
  OAI21X1 U447 ( .A(n1367), .B(n413), .C(n97), .Y(n994) );
  AOI22X1 U448 ( .A(n1027), .B(n215), .C(n300), .D(n995), .Y(n996) );
  NAND3X1 U451 ( .A(n725), .B(n411), .C(n1001), .Y(n1000) );
  NAND3X1 U453 ( .A(counter[0]), .B(n958), .C(n984), .Y(n976) );
  NAND3X1 U454 ( .A(n1004), .B(n1489), .C(n412), .Y(n888) );
  AOI21X1 U455 ( .A(counter[2]), .B(counter[3]), .C(n1491), .Y(n1005) );
  OAI21X1 U456 ( .A(n1007), .B(n1493), .C(n1492), .Y(n1004) );
  NAND3X1 U458 ( .A(n482), .B(n715), .C(n262), .Y(n1010) );
  NAND3X1 U461 ( .A(counter[5]), .B(n1491), .C(n1013), .Y(n889) );
  XNOR2X1 U462 ( .A(n1014), .B(counter[3]), .Y(n1013) );
  NAND3X1 U463 ( .A(n1015), .B(counter[5]), .C(n1014), .Y(n883) );
  NAND3X1 U466 ( .A(n278), .B(n1063), .C(n261), .Y(n1017) );
  AOI22X1 U471 ( .A(n300), .B(n995), .C(n1370), .D(n1027), .Y(n1023) );
  NAND3X1 U473 ( .A(counter[0]), .B(n1025), .C(n1164), .Y(n1022) );
  OAI21X1 U474 ( .A(n476), .B(n433), .C(n116), .Y(n1025) );
  NAND3X1 U475 ( .A(n995), .B(counter[5]), .C(n1029), .Y(n1028) );
  NAND3X1 U478 ( .A(n272), .B(n1063), .C(n1200), .Y(n1031) );
  OAI21X1 U483 ( .A(n211), .B(n247), .C(n1067), .Y(n1043) );
  NAND3X1 U486 ( .A(n1046), .B(n1200), .C(n260), .Y(n1042) );
  NAND3X1 U490 ( .A(n305), .B(n301), .C(n259), .Y(n1049) );
  NAND3X1 U493 ( .A(n1026), .B(n1371), .C(n962), .Y(n1020) );
  NAND3X1 U495 ( .A(n1057), .B(n1063), .C(n1365), .Y(n1056) );
  NAND3X1 U497 ( .A(n1026), .B(n1492), .C(n1007), .Y(n884) );
  OAI21X1 U500 ( .A(n484), .B(n1060), .C(n1067), .Y(n1057) );
  OAI21X1 U501 ( .A(n1048), .B(n995), .C(n1026), .Y(n1060) );
  OAI21X1 U504 ( .A(n415), .B(n243), .C(n140), .Y(n1414) );
  AOI22X1 U506 ( .A(n303), .B(n1503), .C(CMD_data_out[3]), .D(n1068), .Y(n1065) );
  OAI21X1 U507 ( .A(n210), .B(n1504), .C(n115), .Y(n1415) );
  NAND3X1 U508 ( .A(n1068), .B(n1062), .C(CMD_data_out[4]), .Y(n1071) );
  AOI21X1 U510 ( .A(CMD_sz[0]), .B(n303), .C(n415), .Y(n1069) );
  NOR3X1 U512 ( .A(n499), .B(reset), .C(n416), .Y(n1073) );
  AOI22X1 U513 ( .A(n1216), .B(n1027), .C(n1207), .D(n1048), .Y(n1076) );
  AOI22X1 U518 ( .A(CMD_data_out[29]), .B(n1084), .C(n801), .D(n1040), .Y(
        n1083) );
  AOI22X1 U519 ( .A(n611), .B(n1038), .C(n1205), .D(CMD_addr[24]), .Y(n1082)
         );
  AOI22X1 U521 ( .A(CMD_data_out[28]), .B(n1084), .C(n800), .D(n1040), .Y(
        n1091) );
  AOI22X1 U522 ( .A(n610), .B(n1038), .C(n1205), .D(CMD_addr[23]), .Y(n1090)
         );
  AOI22X1 U524 ( .A(CMD_data_out[27]), .B(n1084), .C(n799), .D(n1040), .Y(
        n1093) );
  AOI22X1 U525 ( .A(n609), .B(n1038), .C(n1205), .D(CMD_addr[22]), .Y(n1092)
         );
  AOI22X1 U527 ( .A(CMD_data_out[26]), .B(n1084), .C(n798), .D(n1040), .Y(
        n1095) );
  AOI22X1 U528 ( .A(n608), .B(n1038), .C(n1205), .D(CMD_addr[21]), .Y(n1094)
         );
  AOI22X1 U530 ( .A(CMD_data_out[25]), .B(n1084), .C(n797), .D(n1040), .Y(
        n1097) );
  AOI22X1 U531 ( .A(n607), .B(n1038), .C(n1205), .D(CMD_addr[20]), .Y(n1096)
         );
  AOI22X1 U533 ( .A(CMD_data_out[24]), .B(n1084), .C(n796), .D(n1040), .Y(
        n1099) );
  AOI22X1 U534 ( .A(n606), .B(n1038), .C(n1205), .D(CMD_addr[19]), .Y(n1098)
         );
  AOI22X1 U536 ( .A(CMD_data_out[23]), .B(n1084), .C(n795), .D(n1040), .Y(
        n1101) );
  AOI22X1 U537 ( .A(n605), .B(n1038), .C(n1205), .D(CMD_addr[18]), .Y(n1100)
         );
  AOI22X1 U539 ( .A(CMD_data_out[22]), .B(n1084), .C(n794), .D(n1040), .Y(
        n1103) );
  AOI22X1 U540 ( .A(n604), .B(n1038), .C(n1205), .D(CMD_addr[17]), .Y(n1102)
         );
  AOI22X1 U542 ( .A(CMD_data_out[21]), .B(n1084), .C(n793), .D(n1040), .Y(
        n1105) );
  AOI22X1 U543 ( .A(n603), .B(n1038), .C(n1205), .D(CMD_addr[16]), .Y(n1104)
         );
  AOI22X1 U545 ( .A(CMD_data_out[20]), .B(n1084), .C(n792), .D(n1040), .Y(
        n1119) );
  AOI22X1 U546 ( .A(n602), .B(n1038), .C(n1205), .D(CMD_addr[15]), .Y(n1118)
         );
  AOI22X1 U548 ( .A(CMD_data_out[19]), .B(n1084), .C(n791), .D(n1040), .Y(
        n1122) );
  AOI22X1 U549 ( .A(n601), .B(n1038), .C(n1205), .D(CMD_addr[14]), .Y(n1121)
         );
  AOI22X1 U551 ( .A(CMD_data_out[18]), .B(n1084), .C(n790), .D(n1040), .Y(
        n1124) );
  AOI22X1 U552 ( .A(n600), .B(n1038), .C(n1205), .D(CMD_addr[13]), .Y(n1123)
         );
  AOI22X1 U554 ( .A(CMD_data_out[17]), .B(n1084), .C(n789), .D(n1041), .Y(
        n1126) );
  AOI22X1 U555 ( .A(n599), .B(n1038), .C(n1205), .D(CMD_addr[12]), .Y(n1125)
         );
  AOI22X1 U557 ( .A(CMD_data_out[16]), .B(n1084), .C(n788), .D(n1041), .Y(
        n1128) );
  AOI22X1 U558 ( .A(n598), .B(n1086), .C(n1205), .D(CMD_addr[11]), .Y(n1127)
         );
  AOI22X1 U560 ( .A(CMD_data_out[15]), .B(n1084), .C(n787), .D(n1041), .Y(
        n1130) );
  AOI22X1 U561 ( .A(n597), .B(n1086), .C(n1205), .D(CMD_addr[10]), .Y(n1129)
         );
  AOI22X1 U563 ( .A(CMD_data_out[14]), .B(n1084), .C(n786), .D(n1041), .Y(
        n1132) );
  AOI22X1 U564 ( .A(n596), .B(n1086), .C(n1205), .D(CMD_addr[9]), .Y(n1131) );
  AOI22X1 U566 ( .A(CMD_data_out[13]), .B(n1084), .C(n785), .D(n1041), .Y(
        n1134) );
  AOI22X1 U567 ( .A(n595), .B(n1086), .C(n1205), .D(CMD_addr[8]), .Y(n1133) );
  AOI22X1 U569 ( .A(CMD_data_out[12]), .B(n1084), .C(n784), .D(n1041), .Y(
        n1136) );
  AOI22X1 U570 ( .A(n594), .B(n1086), .C(n1205), .D(CMD_addr[7]), .Y(n1135) );
  AOI22X1 U572 ( .A(CMD_data_out[11]), .B(n1084), .C(n783), .D(n1041), .Y(
        n1138) );
  AOI22X1 U573 ( .A(n593), .B(n1086), .C(n1205), .D(CMD_addr[6]), .Y(n1137) );
  AOI22X1 U575 ( .A(CMD_data_out[10]), .B(n1084), .C(n782), .D(n1041), .Y(
        n1140) );
  AOI22X1 U576 ( .A(n592), .B(n1086), .C(n1205), .D(CMD_addr[5]), .Y(n1139) );
  AOI22X1 U578 ( .A(CMD_data_out[9]), .B(n1084), .C(n781), .D(n1041), .Y(n1142) );
  AOI22X1 U579 ( .A(n591), .B(n1086), .C(n1205), .D(CMD_addr[4]), .Y(n1141) );
  AOI22X1 U581 ( .A(CMD_data_out[8]), .B(n1084), .C(n780), .D(n1041), .Y(n1145) );
  AOI22X1 U582 ( .A(n590), .B(n1086), .C(n1205), .D(CMD_addr[3]), .Y(n1143) );
  AOI22X1 U584 ( .A(CMD_data_out[7]), .B(n1084), .C(n779), .D(n1041), .Y(n1149) );
  AOI22X1 U585 ( .A(n589), .B(n1086), .C(n1205), .D(n762), .Y(n1148) );
  AOI22X1 U587 ( .A(CMD_data_out[6]), .B(n1084), .C(n778), .D(n1041), .Y(n1151) );
  AOI22X1 U588 ( .A(n588), .B(n1086), .C(n1205), .D(n760), .Y(n1150) );
  AOI22X1 U590 ( .A(CMD_data_out[5]), .B(n1084), .C(n777), .D(n1085), .Y(n1153) );
  AOI22X1 U591 ( .A(n587), .B(n1086), .C(n1205), .D(n759), .Y(n1152) );
  AOI22X1 U593 ( .A(CMD_data_out[30]), .B(n1084), .C(n802), .D(n1085), .Y(
        n1155) );
  AOI22X1 U596 ( .A(n612), .B(n1086), .C(n1205), .D(CMD_addr[25]), .Y(n1154)
         );
  OAI21X1 U599 ( .A(reset), .B(n245), .C(n722), .Y(n1157) );
  AOI21X1 U600 ( .A(n1048), .B(n209), .C(n298), .Y(n1158) );
  NAND3X1 U603 ( .A(n1026), .B(counter[3]), .C(n1007), .Y(n1002) );
  NAND3X1 U605 ( .A(n958), .B(n1371), .C(n1026), .Y(n975) );
  NAND3X1 U608 ( .A(n206), .B(n1489), .C(counter[4]), .Y(n1052) );
  NAND3X1 U609 ( .A(n205), .B(n455), .C(n258), .Y(n1162) );
  NAND3X1 U611 ( .A(counter[0]), .B(n958), .C(counter[2]), .Y(n1163) );
  OAI21X1 U613 ( .A(n306), .B(n1053), .C(n101), .Y(n1442) );
  NAND3X1 U614 ( .A(n1169), .B(n1063), .C(n306), .Y(n1168) );
  OAI21X1 U616 ( .A(n1474), .B(n306), .C(n100), .Y(n1443) );
  NAND3X1 U617 ( .A(n306), .B(n1063), .C(n1171), .Y(n1170) );
  OAI21X1 U618 ( .A(n1535), .B(n489), .C(n1174), .Y(n1171) );
  NAND3X1 U620 ( .A(n204), .B(n1554), .C(n1068), .Y(n1175) );
  NAND3X1 U621 ( .A(n489), .B(n1174), .C(n252), .Y(n1176) );
  AOI21X1 U622 ( .A(CMD_data_out[31]), .B(n1537), .C(n1169), .Y(n1177) );
  OAI21X1 U624 ( .A(n1470), .B(n432), .C(n431), .Y(n1444) );
  NAND3X1 U625 ( .A(n1468), .B(n1063), .C(n1184), .Y(n1182) );
  NAND3X1 U628 ( .A(ready), .B(n240), .C(n1187), .Y(n1185) );
  OAI21X1 U630 ( .A(n1033), .B(n1477), .C(n324), .Y(n1445) );
  AOI22X1 U633 ( .A(n218), .B(n1195), .C(we_bar), .D(n723), .Y(n1192) );
  NAND3X1 U634 ( .A(n186), .B(n239), .C(n1198), .Y(n1193) );
  NOR3X1 U635 ( .A(n1473), .B(reset), .C(n1081), .Y(n1198) );
  AOI22X1 U639 ( .A(n1061), .B(n214), .C(n1472), .D(n1202), .Y(n1196) );
  OAI21X1 U642 ( .A(n1479), .B(n1033), .C(n333), .Y(n1447) );
  OAI21X1 U644 ( .A(n1033), .B(n1483), .C(n702), .Y(n1448) );
  OAI21X1 U646 ( .A(n1033), .B(n1484), .C(n406), .Y(n1449) );
  OAI21X1 U648 ( .A(n1485), .B(n1033), .C(n308), .Y(n1450) );
  OAI21X1 U651 ( .A(n1487), .B(n1033), .C(n391), .Y(n1451) );
  OAI21X1 U653 ( .A(n1489), .B(n1033), .C(n342), .Y(n1452) );
  OAI21X1 U655 ( .A(n1491), .B(n1033), .C(n352), .Y(n1453) );
  OAI21X1 U657 ( .A(n1492), .B(n1033), .C(n363), .Y(n1454) );
  OAI21X1 U659 ( .A(n1493), .B(n1033), .C(n427), .Y(n1455) );
  OAI21X1 U661 ( .A(n1494), .B(n1033), .C(n375), .Y(n1456) );
  OAI21X1 U663 ( .A(n1159), .B(n1499), .C(n417), .Y(n1457) );
  OAI21X1 U666 ( .A(n1159), .B(n1498), .C(n381), .Y(n1458) );
  OAI21X1 U669 ( .A(n1159), .B(n1497), .C(n366), .Y(n1459) );
  OAI21X1 U672 ( .A(n1475), .B(n1234), .C(n99), .Y(n1460) );
  NAND3X1 U673 ( .A(n203), .B(n1234), .C(n251), .Y(n1223) );
  AOI21X1 U674 ( .A(CMD_data_out[31]), .B(n1046), .C(n722), .Y(n1225) );
  NAND3X1 U675 ( .A(n1536), .B(n1537), .C(n1535), .Y(n1224) );
  OAI21X1 U676 ( .A(n1054), .B(n1234), .C(n96), .Y(n1461) );
  AOI22X1 U677 ( .A(n1209), .B(n863), .C(n1159), .D(n1169), .Y(n1227) );
  OAI21X1 U678 ( .A(n460), .B(n1535), .C(n139), .Y(n1169) );
  OAI21X1 U682 ( .A(refresh_counter[12]), .B(n1470), .C(n681), .Y(n863) );
  NAND3X1 U685 ( .A(n1231), .B(n238), .C(n257), .Y(n1462) );
  NAND3X1 U687 ( .A(n1234), .B(n1535), .C(n250), .Y(n1232) );
  AOI21X1 U688 ( .A(n460), .B(n489), .C(n722), .Y(n1235) );
  NOR3X1 U690 ( .A(state[0]), .B(state[2]), .C(n1054), .Y(n1068) );
  OAI21X1 U696 ( .A(refresh_counter[12]), .B(n1470), .C(n1209), .Y(n1231) );
  NAND3X1 U698 ( .A(n1234), .B(n1063), .C(n1187), .Y(n1236) );
  OAI21X1 U702 ( .A(n711), .B(n1468), .C(n463), .Y(n1463) );
  AOI21X1 U708 ( .A(n1473), .B(n1373), .C(reset), .Y(n1238) );
  NOR3X1 U709 ( .A(n1487), .B(n458), .C(n408), .Y(n1373) );
  OAI21X1 U712 ( .A(n1371), .B(n1033), .C(n315), .Y(n1464) );
  NAND3X1 U716 ( .A(n494), .B(n456), .C(n1244), .Y(n1188) );
  NOR3X1 U717 ( .A(n1472), .B(reset), .C(n1187), .Y(n1244) );
  NOR3X1 U718 ( .A(state[1]), .B(state[2]), .C(state[0]), .Y(n1187) );
  NAND3X1 U720 ( .A(n1054), .B(n1475), .C(state[0]), .Y(n833) );
  NAND3X1 U721 ( .A(state[0]), .B(n1475), .C(state[1]), .Y(n1242) );
  NAND3X1 U726 ( .A(state[2]), .B(n1054), .C(state[0]), .Y(n1080) );
  OAI21X1 U729 ( .A(n1147), .B(reset), .C(n1195), .Y(n1246) );
  OAI21X1 U732 ( .A(n1146), .B(reset), .C(n1195), .Y(n1248) );
  NOR3X1 U736 ( .A(n365), .B(n435), .C(n462), .Y(n890) );
  AOI21X1 U737 ( .A(n434), .B(n1363), .C(n462), .Y(n881) );
  NAND3X1 U752 ( .A(counter[4]), .B(n1493), .C(n1253), .Y(n1249) );
  NOR3X1 U753 ( .A(n378), .B(n435), .C(n462), .Y(n648) );
  AOI21X1 U767 ( .A(n1504), .B(n1503), .C(n1474), .Y(n1079) );
  NAND3X1 U773 ( .A(counter[2]), .B(n1491), .C(n1253), .Y(n1254) );
  NOR3X1 U774 ( .A(n484), .B(n1371), .C(n1489), .Y(n1253) );
  AOI21X1 U775 ( .A(n287), .B(n208), .C(n458), .Y(n350) );
  NAND3X1 U776 ( .A(n1360), .B(n1479), .C(n1257), .Y(n1240) );
  NOR3X1 U777 ( .A(counter[2]), .B(counter[7]), .C(counter[5]), .Y(n1257) );
  NAND3X1 U779 ( .A(n1491), .B(n1487), .C(n1059), .Y(n1256) );
  NAND3X1 U780 ( .A(n1491), .B(n1487), .C(n958), .Y(n866) );
  NOR3X1 U781 ( .A(n710), .B(n479), .C(n1479), .Y(n284) );
  NAND3X1 U783 ( .A(n1484), .B(n1483), .C(n1260), .Y(n1258) );
  NAND3X1 U788 ( .A(n1482), .B(n1059), .C(counter[5]), .Y(n844) );
  OAI21X1 U792 ( .A(counter[10]), .B(n244), .C(n138), .Y(n1202) );
  NAND3X1 U795 ( .A(counter[4]), .B(counter[2]), .C(n960), .Y(n1265) );
  AOI21X1 U796 ( .A(n1266), .B(n1487), .C(n1486), .Y(n1263) );
  NAND3X1 U798 ( .A(counter[7]), .B(n1494), .C(n1268), .Y(n1259) );
  OAI21X1 U801 ( .A(counter[7]), .B(n242), .C(n98), .Y(n1266) );
  NAND3X1 U802 ( .A(n1164), .B(counter[7]), .C(n1490), .Y(n1271) );
  AOI22X1 U806 ( .A(n961), .B(n962), .C(n1488), .D(counter[1]), .Y(n1270) );
  NAND3X1 U807 ( .A(n960), .B(n1494), .C(n1488), .Y(n832) );
  OAI21X1 U808 ( .A(ATOMIC_cmd), .B(n1553), .C(n317), .Y(n1391) );
  OAI21X1 U811 ( .A(ATOMIC_cmd), .B(n1552), .C(n326), .Y(n1390) );
  OAI21X1 U814 ( .A(ATOMIC_cmd), .B(n1551), .C(n355), .Y(n1389) );
  OAI21X1 U817 ( .A(ATOMIC_cmd), .B(n1550), .C(n367), .Y(n1388) );
  OAI21X1 U820 ( .A(ATOMIC_cmd), .B(n1549), .C(n383), .Y(n1387) );
  OAI21X1 U823 ( .A(ATOMIC_cmd), .B(n1548), .C(n398), .Y(n1386) );
  OAI21X1 U826 ( .A(ATOMIC_cmd), .B(n1547), .C(n335), .Y(n1385) );
  OAI21X1 U829 ( .A(ATOMIC_cmd), .B(n1546), .C(n344), .Y(n1384) );
  OAI21X1 U832 ( .A(ATOMIC_cmd), .B(n1545), .C(n356), .Y(n1383) );
  OAI21X1 U835 ( .A(ATOMIC_cmd), .B(n1544), .C(n368), .Y(n1382) );
  OAI21X1 U838 ( .A(ATOMIC_cmd), .B(n1543), .C(n384), .Y(n1381) );
  OAI21X1 U841 ( .A(ATOMIC_cmd), .B(n1542), .C(n399), .Y(n1380) );
  OAI21X1 U844 ( .A(ATOMIC_cmd), .B(n1541), .C(n420), .Y(n1379) );
  OAI21X1 U847 ( .A(ATOMIC_cmd), .B(n1540), .C(n437), .Y(n1378) );
  OAI21X1 U850 ( .A(ATOMIC_cmd), .B(n1539), .C(n465), .Y(n1377) );
  OAI21X1 U853 ( .A(ATOMIC_cmd), .B(n1538), .C(n673), .Y(n1376) );
  AOI21X1 U856 ( .A(n434), .B(n1362), .C(n462), .Y(n1088) );
  NOR3X1 U858 ( .A(n290), .B(n462), .C(n394), .Y(n1087) );
  NAND3X1 U859 ( .A(counter[4]), .B(n1493), .C(counter[5]), .Y(n1273) );
  NAND3X1 U860 ( .A(n960), .B(n1477), .C(n1291), .Y(n1250) );
  NOR3X1 U865 ( .A(counter[6]), .B(counter[7]), .C(counter[10]), .Y(n960) );
  NAND3X1 U869 ( .A(n396), .B(n1363), .C(n724), .Y(n1064) );
  OAI21X1 U871 ( .A(counter[0]), .B(n395), .C(n461), .Y(n835) );
  NAND3X1 U872 ( .A(n1015), .B(n1161), .C(n1007), .Y(n829) );
  NAND3X1 U873 ( .A(n1007), .B(n1492), .C(n984), .Y(n830) );
  OAI21X1 U876 ( .A(counter[0]), .B(n395), .C(n434), .Y(n834) );
  AOI21X1 U880 ( .A(counter[1]), .B(n1488), .C(n1293), .Y(n1292) );
  NAND3X1 U885 ( .A(n1493), .B(n1489), .C(n1015), .Y(n1294) );
  NAND3X1 U890 ( .A(n958), .B(n1371), .C(n984), .Y(n999) );
  NOR3X1 U891 ( .A(counter[2]), .B(counter[5]), .C(n1491), .Y(n984) );
  ddr3_ring_buffer8 ring_buffer ( .dout(RETURN_data), .listen(listen), 
        .strobe(DQS_in), .readPtr(read_pointer), .din(DQ_in), .reset(reset) );
  Processing_logic_DW01_add_0 add_663 ( .A(RETURN_data), .B(DATA_data_out), 
        .CI(1'b0), .SUM({n1325, n1324, n1323, n1322, n1321, n1320, n1319, 
        n1318, n1317, n1316, n1315, n1314, n1313, n1312, n1311, n1310}), .CO()
         );
  Processing_logic_DW01_add_2 add_526 ( .A({CMD_addr, n762, n760, n759}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 
        1'b0, 1'b0}), .CI(1'b0), .SUM({n802, n801, n800, n799, n798, n797, 
        n796, n795, n794, n793, n792, n791, n790, n789, n788, n787, n786, n785, 
        n784, n783, n782, n781, n780, n779, n778, n777}), .CO() );
  Processing_logic_DW01_inc_0 add_185 ( .A(refresh_counter), .SUM({n114, n113, 
        n112, n111, n110, n109, n108, n107, n106, n105, n104, n103, n102}) );
  Processing_logic_DW01_inc_1 r474 ( .A({CMD_addr, n762, n760, n759}), .SUM({
        n612, n611, n610, n609, n608, n607, n606, n605, n604, n603, n602, n601, 
        n600, n599, n598, n597, n596, n595, n594, n593, n592, n591, n590, n589, 
        n588, n587}) );
  Processing_logic_DW01_inc_2 r473 ( .A(counter), .SUM({n163, n162, n161, n160, 
        n159, n158, n157, n156, n155, n154, n153, n152}) );
  AND2X1 U4 ( .A(n153), .B(n728), .Y(n629) );
  AND2X1 U7 ( .A(n154), .B(n728), .Y(n630) );
  AND2X1 U11 ( .A(n155), .B(n728), .Y(n631) );
  AND2X1 U15 ( .A(n156), .B(n728), .Y(n632) );
  AND2X1 U22 ( .A(n157), .B(n728), .Y(n633) );
  AND2X1 U24 ( .A(n158), .B(n728), .Y(n634) );
  AND2X1 U28 ( .A(n160), .B(n728), .Y(n636) );
  AND2X1 U29 ( .A(n161), .B(n728), .Y(n637) );
  AND2X1 U35 ( .A(n162), .B(n728), .Y(n638) );
  AND2X1 U39 ( .A(n163), .B(n728), .Y(n639) );
  AND2X1 U45 ( .A(n152), .B(n728), .Y(n628) );
  AND2X1 U49 ( .A(n302), .B(n307), .Y(n926) );
  AND2X1 U55 ( .A(n304), .B(n307), .Y(n927) );
  OR2X1 U59 ( .A(n285), .B(n433), .Y(n895) );
  AND2X1 U65 ( .A(state[1]), .B(n720), .Y(n1061) );
  AND2X1 U69 ( .A(n62), .B(n716), .Y(n719) );
  AND2X1 U75 ( .A(counter[0]), .B(n720), .Y(n726) );
  OR2X1 U79 ( .A(n184), .B(n185), .Y(n941) );
  AND2X1 U85 ( .A(n159), .B(n728), .Y(n635) );
  AND2X1 U89 ( .A(n159), .B(n498), .Y(n876) );
  AND2X1 U95 ( .A(n414), .B(n276), .Y(n275) );
  OR2X1 U99 ( .A(n816), .B(n494), .Y(n818) );
  OR2X1 U105 ( .A(n414), .B(n481), .Y(n824) );
  AND2X1 U109 ( .A(n153), .B(n498), .Y(n870) );
  AND2X1 U115 ( .A(n154), .B(n498), .Y(n871) );
  AND2X1 U119 ( .A(n155), .B(n498), .Y(n872) );
  AND2X1 U125 ( .A(n156), .B(n498), .Y(n873) );
  AND2X1 U129 ( .A(n157), .B(n498), .Y(n874) );
  AND2X1 U135 ( .A(n158), .B(n498), .Y(n875) );
  AND2X1 U139 ( .A(n160), .B(n498), .Y(n877) );
  AND2X1 U145 ( .A(n161), .B(n498), .Y(n878) );
  AND2X1 U149 ( .A(n162), .B(n498), .Y(n879) );
  AND2X1 U155 ( .A(n163), .B(n498), .Y(n880) );
  OR2X1 U159 ( .A(n460), .B(CMD_data_out[31]), .Y(n1174) );
  AND2X1 U163 ( .A(n1063), .B(n93), .Y(n1166) );
  AND2X1 U164 ( .A(n1067), .B(n92), .Y(n1181) );
  AND2X1 U166 ( .A(n152), .B(n498), .Y(n869) );
  AND2X1 U170 ( .A(n61), .B(n91), .Y(n506) );
  AND2X1 U172 ( .A(n60), .B(n90), .Y(n518) );
  AND2X1 U173 ( .A(n59), .B(n89), .Y(n528) );
  AND2X1 U175 ( .A(n58), .B(n88), .Y(n538) );
  AND2X1 U177 ( .A(n57), .B(n87), .Y(n548) );
  AND2X1 U179 ( .A(n56), .B(n86), .Y(n558) );
  AND2X1 U181 ( .A(n55), .B(n85), .Y(n568) );
  AND2X1 U183 ( .A(n54), .B(n84), .Y(n578) );
  AND2X1 U187 ( .A(n53), .B(n83), .Y(n614) );
  AND2X1 U188 ( .A(n52), .B(n82), .Y(n624) );
  AND2X1 U190 ( .A(n51), .B(n81), .Y(n646) );
  AND2X1 U192 ( .A(n50), .B(n80), .Y(n657) );
  AND2X1 U197 ( .A(n49), .B(n79), .Y(n667) );
  AND2X1 U198 ( .A(n48), .B(n78), .Y(n677) );
  AND2X1 U199 ( .A(n698), .B(n693), .Y(n1417) );
  AND2X1 U201 ( .A(n443), .B(n442), .Y(n1418) );
  AND2X1 U202 ( .A(n426), .B(n425), .Y(n1419) );
  AND2X1 U204 ( .A(n405), .B(n404), .Y(n1420) );
  AND2X1 U206 ( .A(n390), .B(n389), .Y(n1421) );
  AND2X1 U207 ( .A(n374), .B(n373), .Y(n1422) );
  AND2X1 U209 ( .A(n362), .B(n361), .Y(n1423) );
  AND2X1 U211 ( .A(n351), .B(n349), .Y(n1424) );
  AND2X1 U213 ( .A(n341), .B(n340), .Y(n1425) );
  AND2X1 U214 ( .A(n332), .B(n331), .Y(n1426) );
  AND2X1 U216 ( .A(n323), .B(n322), .Y(n1427) );
  AND2X1 U217 ( .A(n313), .B(n314), .Y(n1428) );
  AND2X1 U219 ( .A(n422), .B(n423), .Y(n1429) );
  AND2X1 U220 ( .A(n401), .B(n402), .Y(n1430) );
  AND2X1 U222 ( .A(n386), .B(n387), .Y(n1431) );
  AND2X1 U223 ( .A(n370), .B(n371), .Y(n1432) );
  AND2X1 U225 ( .A(n358), .B(n359), .Y(n1433) );
  AND2X1 U226 ( .A(n346), .B(n347), .Y(n1434) );
  AND2X1 U228 ( .A(n337), .B(n338), .Y(n1435) );
  AND2X1 U229 ( .A(n328), .B(n329), .Y(n1436) );
  AND2X1 U231 ( .A(n469), .B(n470), .Y(n1437) );
  AND2X1 U232 ( .A(n319), .B(n320), .Y(n1438) );
  AND2X1 U234 ( .A(n310), .B(n311), .Y(n1439) );
  AND2X1 U235 ( .A(n447), .B(n448), .Y(n1440) );
  AND2X1 U237 ( .A(n473), .B(n472), .Y(n1416) );
  AND2X1 U238 ( .A(n686), .B(n685), .Y(n1441) );
  AND2X1 U240 ( .A(n440), .B(n439), .Y(n1413) );
  AND2X1 U241 ( .A(n467), .B(n1246), .Y(n1465) );
  AND2X1 U243 ( .A(n445), .B(n1248), .Y(n1466) );
  AND2X1 U244 ( .A(n816), .B(n94), .Y(n930) );
  AND2X1 U246 ( .A(n1067), .B(n95), .Y(n822) );
  AND2X1 U247 ( .A(n267), .B(n268), .Y(n831) );
  AND2X1 U249 ( .A(n47), .B(n1446), .Y(n973) );
  AND2X1 U250 ( .A(n430), .B(n1058), .Y(n860) );
  AND2X1 U252 ( .A(n1480), .B(n379), .Y(n276) );
  XOR2X1 U253 ( .A(counter[3]), .B(n762), .Y(n1) );
  BUFX2 U255 ( .A(n1326), .Y(n2) );
  BUFX2 U256 ( .A(n1309), .Y(n3) );
  BUFX2 U258 ( .A(n1308), .Y(n4) );
  BUFX2 U259 ( .A(n1307), .Y(n5) );
  BUFX2 U261 ( .A(n1306), .Y(n6) );
  BUFX2 U262 ( .A(n1305), .Y(n7) );
  BUFX2 U264 ( .A(n1304), .Y(n8) );
  BUFX2 U265 ( .A(n1303), .Y(n9) );
  BUFX2 U267 ( .A(n1302), .Y(n10) );
  BUFX2 U269 ( .A(n1301), .Y(n11) );
  BUFX2 U271 ( .A(n1300), .Y(n12) );
  BUFX2 U272 ( .A(n1299), .Y(n13) );
  BUFX2 U274 ( .A(n1298), .Y(n14) );
  BUFX2 U276 ( .A(n1297), .Y(n15) );
  BUFX2 U277 ( .A(n1296), .Y(n16) );
  BUFX2 U278 ( .A(n1295), .Y(n17) );
  BUFX2 U280 ( .A(n1192), .Y(n18) );
  BUFX2 U281 ( .A(n1023), .Y(n19) );
  BUFX2 U286 ( .A(n859), .Y(n20) );
  BUFX2 U287 ( .A(n858), .Y(n21) );
  BUFX2 U288 ( .A(n857), .Y(n22) );
  BUFX2 U289 ( .A(n856), .Y(n23) );
  BUFX2 U292 ( .A(n855), .Y(n24) );
  BUFX2 U294 ( .A(n854), .Y(n25) );
  BUFX2 U295 ( .A(n853), .Y(n26) );
  BUFX2 U297 ( .A(n852), .Y(n27) );
  BUFX2 U299 ( .A(n851), .Y(n28) );
  BUFX2 U301 ( .A(n850), .Y(n29) );
  BUFX2 U303 ( .A(n849), .Y(n30) );
  BUFX2 U305 ( .A(n846), .Y(n31) );
  AND2X1 U307 ( .A(n430), .B(n711), .Y(n847) );
  BUFX2 U309 ( .A(n819), .Y(n32) );
  BUFX2 U311 ( .A(n1294), .Y(n33) );
  BUFX2 U313 ( .A(n1265), .Y(n34) );
  BUFX2 U315 ( .A(n1236), .Y(n35) );
  BUFX2 U317 ( .A(n1042), .Y(n36) );
  BUFX2 U319 ( .A(n1022), .Y(n37) );
  BUFX2 U320 ( .A(n1010), .Y(n38) );
  BUFX2 U322 ( .A(n1000), .Y(n39) );
  AND2X1 U324 ( .A(n285), .B(n299), .Y(n1001) );
  BUFX2 U329 ( .A(n956), .Y(n40) );
  BUFX2 U330 ( .A(n891), .Y(n41) );
  BUFX2 U334 ( .A(n892), .Y(n42) );
  BUFX2 U335 ( .A(n718), .Y(n43) );
  BUFX2 U336 ( .A(n695), .Y(n44) );
  OR2X1 U337 ( .A(n1034), .B(n277), .Y(n273) );
  INVX1 U339 ( .A(n273), .Y(n45) );
  OR2X1 U343 ( .A(n1043), .B(n274), .Y(n277) );
  OR2X1 U345 ( .A(n281), .B(n282), .Y(n279) );
  INVX1 U346 ( .A(n279), .Y(n46) );
  OR2X1 U347 ( .A(n280), .B(reset), .Y(n282) );
  OR2X1 U349 ( .A(n295), .B(n297), .Y(n292) );
  OR2X1 U354 ( .A(n293), .B(n294), .Y(n297) );
  AND2X1 U355 ( .A(n1048), .B(n148), .Y(n1034) );
  BUFX2 U356 ( .A(n978), .Y(n47) );
  BUFX2 U357 ( .A(n678), .Y(n48) );
  BUFX2 U358 ( .A(n668), .Y(n49) );
  BUFX2 U360 ( .A(n658), .Y(n50) );
  BUFX2 U361 ( .A(n647), .Y(n51) );
  BUFX2 U363 ( .A(n625), .Y(n52) );
  BUFX2 U364 ( .A(n615), .Y(n53) );
  BUFX2 U366 ( .A(n579), .Y(n54) );
  BUFX2 U367 ( .A(n569), .Y(n55) );
  BUFX2 U369 ( .A(n559), .Y(n56) );
  BUFX2 U370 ( .A(n549), .Y(n57) );
  BUFX2 U371 ( .A(n539), .Y(n58) );
  BUFX2 U372 ( .A(n529), .Y(n59) );
  BUFX2 U373 ( .A(n519), .Y(n60) );
  BUFX2 U375 ( .A(n507), .Y(n61) );
  BUFX2 U378 ( .A(n721), .Y(n62) );
  BUFX2 U379 ( .A(n1462), .Y(n63) );
  AND2X1 U381 ( .A(n181), .B(n149), .Y(n1412) );
  INVX1 U382 ( .A(n1412), .Y(n64) );
  AND2X1 U384 ( .A(n182), .B(n150), .Y(n1411) );
  INVX1 U385 ( .A(n1411), .Y(n65) );
  AND2X1 U387 ( .A(n183), .B(n151), .Y(n1408) );
  INVX1 U389 ( .A(n1408), .Y(n66) );
  AND2X1 U390 ( .A(n170), .B(n164), .Y(n1406) );
  INVX1 U392 ( .A(n1406), .Y(n67) );
  AND2X1 U395 ( .A(n171), .B(n143), .Y(n1405) );
  INVX1 U398 ( .A(n1405), .Y(n68) );
  AND2X1 U399 ( .A(n172), .B(n144), .Y(n1404) );
  INVX1 U402 ( .A(n1404), .Y(n69) );
  AND2X1 U403 ( .A(n173), .B(n145), .Y(n1403) );
  INVX1 U404 ( .A(n1403), .Y(n70) );
  AND2X1 U405 ( .A(n174), .B(n146), .Y(n1402) );
  INVX1 U407 ( .A(n1402), .Y(n71) );
  AND2X1 U408 ( .A(n175), .B(n165), .Y(n1401) );
  INVX1 U409 ( .A(n1401), .Y(n72) );
  AND2X1 U411 ( .A(n176), .B(n166), .Y(n1400) );
  INVX1 U412 ( .A(n1400), .Y(n73) );
  AND2X1 U414 ( .A(n177), .B(n167), .Y(n1399) );
  INVX1 U416 ( .A(n1399), .Y(n74) );
  AND2X1 U421 ( .A(n178), .B(n147), .Y(n1398) );
  INVX1 U424 ( .A(n1398), .Y(n75) );
  AND2X1 U425 ( .A(n179), .B(n168), .Y(n1397) );
  INVX1 U427 ( .A(n1397), .Y(n76) );
  AND2X1 U428 ( .A(n180), .B(n169), .Y(n1356) );
  INVX1 U429 ( .A(n1356), .Y(n77) );
  BUFX2 U431 ( .A(n679), .Y(n78) );
  BUFX2 U432 ( .A(n669), .Y(n79) );
  BUFX2 U433 ( .A(n659), .Y(n80) );
  BUFX2 U434 ( .A(n649), .Y(n81) );
  BUFX2 U438 ( .A(n626), .Y(n82) );
  BUFX2 U441 ( .A(n616), .Y(n83) );
  BUFX2 U444 ( .A(n580), .Y(n84) );
  BUFX2 U445 ( .A(n570), .Y(n85) );
  BUFX2 U446 ( .A(n560), .Y(n86) );
  BUFX2 U449 ( .A(n550), .Y(n87) );
  BUFX2 U450 ( .A(n540), .Y(n88) );
  BUFX2 U452 ( .A(n530), .Y(n89) );
  BUFX2 U457 ( .A(n520), .Y(n90) );
  BUFX2 U459 ( .A(n508), .Y(n91) );
  BUFX2 U460 ( .A(n1185), .Y(n92) );
  BUFX2 U464 ( .A(n1175), .Y(n93) );
  BUFX2 U465 ( .A(n954), .Y(n94) );
  BUFX2 U467 ( .A(n836), .Y(n95) );
  BUFX2 U468 ( .A(n1227), .Y(n96) );
  BUFX2 U469 ( .A(n996), .Y(n97) );
  BUFX2 U470 ( .A(n1271), .Y(n98) );
  BUFX2 U472 ( .A(n1223), .Y(n99) );
  BUFX2 U476 ( .A(n1170), .Y(n100) );
  BUFX2 U477 ( .A(n1168), .Y(n101) );
  BUFX2 U479 ( .A(n1071), .Y(n115) );
  BUFX2 U480 ( .A(n1028), .Y(n116) );
  BUFX2 U481 ( .A(n991), .Y(n117) );
  BUFX2 U482 ( .A(n988), .Y(n118) );
  BUFX2 U484 ( .A(n982), .Y(n119) );
  BUFX2 U485 ( .A(n868), .Y(n120) );
  BUFX2 U487 ( .A(n717), .Y(n121) );
  BUFX2 U488 ( .A(n700), .Y(n122) );
  BUFX2 U489 ( .A(n684), .Y(n123) );
  BUFX2 U491 ( .A(n674), .Y(n124) );
  BUFX2 U492 ( .A(n664), .Y(n125) );
  BUFX2 U494 ( .A(n654), .Y(n126) );
  BUFX2 U496 ( .A(n643), .Y(n127) );
  BUFX2 U498 ( .A(n621), .Y(n128) );
  BUFX2 U499 ( .A(n585), .Y(n129) );
  BUFX2 U502 ( .A(n575), .Y(n130) );
  BUFX2 U503 ( .A(n565), .Y(n131) );
  BUFX2 U505 ( .A(n555), .Y(n132) );
  BUFX2 U509 ( .A(n545), .Y(n133) );
  BUFX2 U511 ( .A(n535), .Y(n134) );
  BUFX2 U514 ( .A(n525), .Y(n135) );
  BUFX2 U515 ( .A(n514), .Y(n136) );
  BUFX2 U516 ( .A(n497), .Y(n137) );
  AND2X1 U517 ( .A(n1482), .B(n958), .Y(n1264) );
  INVX1 U520 ( .A(n1264), .Y(n138) );
  AND2X1 U523 ( .A(n1046), .B(n1535), .Y(n1229) );
  INVX1 U526 ( .A(n1229), .Y(n139) );
  AND2X1 U529 ( .A(CMD_sz[0]), .B(n415), .Y(n1066) );
  INVX1 U532 ( .A(n1066), .Y(n140) );
  AND2X1 U535 ( .A(RETURN_data[1]), .B(n1495), .Y(n694) );
  INVX1 U538 ( .A(n694), .Y(n141) );
  AND2X1 U541 ( .A(RETURN_data[7]), .B(n1024), .Y(n491) );
  INVX1 U544 ( .A(n491), .Y(n142) );
  BUFX2 U547 ( .A(n949), .Y(n143) );
  BUFX2 U550 ( .A(n946), .Y(n144) );
  BUFX2 U553 ( .A(n943), .Y(n145) );
  BUFX2 U556 ( .A(n939), .Y(n146) );
  BUFX2 U559 ( .A(n929), .Y(n147) );
  BUFX2 U562 ( .A(n1049), .Y(n148) );
  BUFX2 U565 ( .A(n1031), .Y(n149) );
  BUFX2 U568 ( .A(n1017), .Y(n150) );
  BUFX2 U571 ( .A(n972), .Y(n151) );
  AND2X1 U574 ( .A(A[0]), .B(n930), .Y(n953) );
  INVX1 U577 ( .A(n953), .Y(n164) );
  AND2X1 U580 ( .A(A[5]), .B(n930), .Y(n937) );
  INVX1 U583 ( .A(n937), .Y(n165) );
  AND2X1 U586 ( .A(A[6]), .B(n930), .Y(n935) );
  INVX1 U589 ( .A(n935), .Y(n166) );
  AND2X1 U592 ( .A(A[7]), .B(n930), .Y(n933) );
  INVX1 U594 ( .A(n933), .Y(n167) );
  AND2X1 U595 ( .A(A[9]), .B(n930), .Y(n924) );
  INVX1 U597 ( .A(n924), .Y(n168) );
  AND2X1 U598 ( .A(BA[0]), .B(n816), .Y(n813) );
  INVX1 U601 ( .A(n813), .Y(n169) );
  BUFX2 U602 ( .A(n952), .Y(n170) );
  BUFX2 U604 ( .A(n948), .Y(n171) );
  BUFX2 U606 ( .A(n945), .Y(n172) );
  BUFX2 U607 ( .A(n942), .Y(n173) );
  BUFX2 U610 ( .A(n938), .Y(n174) );
  BUFX2 U612 ( .A(n936), .Y(n175) );
  BUFX2 U615 ( .A(n934), .Y(n176) );
  BUFX2 U619 ( .A(n932), .Y(n177) );
  BUFX2 U623 ( .A(n928), .Y(n178) );
  BUFX2 U626 ( .A(n923), .Y(n179) );
  BUFX2 U627 ( .A(n812), .Y(n180) );
  AND2X1 U629 ( .A(RETURN_put), .B(n45), .Y(n1030) );
  INVX1 U631 ( .A(n1030), .Y(n181) );
  AND2X1 U632 ( .A(ts_con), .B(n46), .Y(n1016) );
  INVX1 U636 ( .A(n1016), .Y(n182) );
  AND2X1 U637 ( .A(DATA_get), .B(n973), .Y(n971) );
  INVX1 U638 ( .A(n971), .Y(n183) );
  BUFX2 U640 ( .A(n965), .Y(n184) );
  BUFX2 U641 ( .A(n966), .Y(n185) );
  BUFX2 U643 ( .A(n1196), .Y(n186) );
  BUFX2 U645 ( .A(n689), .Y(n187) );
  BUFX2 U647 ( .A(n675), .Y(n188) );
  BUFX2 U649 ( .A(n665), .Y(n189) );
  BUFX2 U650 ( .A(n655), .Y(n190) );
  BUFX2 U652 ( .A(n644), .Y(n191) );
  BUFX2 U654 ( .A(n622), .Y(n192) );
  BUFX2 U656 ( .A(n586), .Y(n193) );
  BUFX2 U658 ( .A(n576), .Y(n194) );
  BUFX2 U660 ( .A(n566), .Y(n195) );
  BUFX2 U662 ( .A(n556), .Y(n196) );
  BUFX2 U664 ( .A(n546), .Y(n197) );
  BUFX2 U665 ( .A(n536), .Y(n198) );
  BUFX2 U667 ( .A(n526), .Y(n199) );
  BUFX2 U668 ( .A(n516), .Y(n200) );
  BUFX2 U670 ( .A(n504), .Y(n201) );
  BUFX2 U671 ( .A(n485), .Y(n202) );
  BUFX2 U679 ( .A(n1224), .Y(n203) );
  BUFX2 U680 ( .A(n1176), .Y(n204) );
  BUFX2 U681 ( .A(n1163), .Y(n205) );
  BUFX2 U683 ( .A(n1162), .Y(n206) );
  INVX1 U684 ( .A(n719), .Y(n207) );
  BUFX2 U686 ( .A(n1256), .Y(n208) );
  AND2X1 U689 ( .A(n271), .B(n305), .Y(n1160) );
  INVX1 U691 ( .A(n1160), .Y(n209) );
  BUFX2 U692 ( .A(n1069), .Y(n210) );
  AND2X1 U693 ( .A(counter[0]), .B(n958), .Y(n1044) );
  INVX1 U694 ( .A(n1044), .Y(n211) );
  OR2X1 U695 ( .A(n998), .B(n828), .Y(n841) );
  INVX1 U697 ( .A(n841), .Y(n212) );
  BUFX2 U699 ( .A(n821), .Y(n213) );
  AND2X1 U700 ( .A(n461), .B(n409), .Y(n1201) );
  INVX1 U701 ( .A(n1201), .Y(n214) );
  AND2X1 U703 ( .A(n1364), .B(n724), .Y(n997) );
  INVX1 U704 ( .A(n997), .Y(n215) );
  BUFX2 U705 ( .A(n1088), .Y(n216) );
  BUFX2 U706 ( .A(n350), .Y(n217) );
  BUFX2 U707 ( .A(n1193), .Y(n218) );
  BUFX2 U710 ( .A(n840), .Y(n219) );
  AND2X1 U711 ( .A(n1478), .B(n941), .Y(n940) );
  INVX1 U713 ( .A(n940), .Y(n220) );
  AND2X1 U714 ( .A(n411), .B(n715), .Y(n886) );
  INVX1 U715 ( .A(n886), .Y(n221) );
  BUFX2 U719 ( .A(n690), .Y(n222) );
  BUFX2 U722 ( .A(n676), .Y(n223) );
  BUFX2 U723 ( .A(n666), .Y(n224) );
  BUFX2 U724 ( .A(n656), .Y(n225) );
  BUFX2 U725 ( .A(n645), .Y(n226) );
  BUFX2 U727 ( .A(n623), .Y(n227) );
  BUFX2 U728 ( .A(n613), .Y(n228) );
  BUFX2 U730 ( .A(n577), .Y(n229) );
  BUFX2 U731 ( .A(n567), .Y(n230) );
  BUFX2 U733 ( .A(n557), .Y(n231) );
  BUFX2 U734 ( .A(n547), .Y(n232) );
  BUFX2 U735 ( .A(n537), .Y(n233) );
  BUFX2 U738 ( .A(n527), .Y(n234) );
  BUFX2 U739 ( .A(n517), .Y(n235) );
  BUFX2 U740 ( .A(n505), .Y(n236) );
  BUFX2 U741 ( .A(n486), .Y(n237) );
  BUFX2 U742 ( .A(n1232), .Y(n238) );
  AND2X1 U743 ( .A(n266), .B(n834), .Y(n1197) );
  INVX1 U744 ( .A(n1197), .Y(n239) );
  AND2X1 U745 ( .A(CMD_empty), .B(n1470), .Y(n1186) );
  INVX1 U746 ( .A(n1186), .Y(n240) );
  AND2X1 U747 ( .A(n302), .B(n1476), .Y(n838) );
  INVX1 U748 ( .A(n838), .Y(n241) );
  BUFX2 U749 ( .A(n1270), .Y(n242) );
  BUFX2 U750 ( .A(n1065), .Y(n243) );
  BUFX2 U751 ( .A(n1263), .Y(n244) );
  BUFX2 U754 ( .A(n1158), .Y(n245) );
  BUFX2 U755 ( .A(n903), .Y(n246) );
  AND2X1 U756 ( .A(n995), .B(n1026), .Y(n1045) );
  INVX1 U757 ( .A(n1045), .Y(n247) );
  BUFX2 U758 ( .A(n885), .Y(n248) );
  BUFX2 U759 ( .A(n839), .Y(n249) );
  BUFX2 U760 ( .A(n1235), .Y(n250) );
  BUFX2 U761 ( .A(n1225), .Y(n251) );
  BUFX2 U762 ( .A(n1177), .Y(n252) );
  BUFX2 U763 ( .A(n882), .Y(n253) );
  BUFX2 U764 ( .A(n825), .Y(n254) );
  BUFX2 U765 ( .A(n691), .Y(n255) );
  BUFX2 U766 ( .A(n487), .Y(n256) );
  AND2X1 U768 ( .A(n475), .B(state[0]), .Y(n1233) );
  INVX1 U769 ( .A(n1233), .Y(n257) );
  AND2X1 U770 ( .A(counter[3]), .B(n1493), .Y(n1165) );
  INVX1 U771 ( .A(n1165), .Y(n258) );
  AND2X1 U772 ( .A(n1467), .B(n1474), .Y(n1050) );
  INVX1 U778 ( .A(n1050), .Y(n259) );
  OR2X1 U782 ( .A(n413), .B(CMD_data_out[31]), .Y(n1047) );
  INVX1 U784 ( .A(n1047), .Y(n260) );
  AND2X1 U785 ( .A(n724), .B(n301), .Y(n1019) );
  INVX1 U786 ( .A(n1019), .Y(n261) );
  AND2X1 U787 ( .A(n1012), .B(n1026), .Y(n1011) );
  INVX1 U789 ( .A(n1011), .Y(n262) );
  AND2X1 U790 ( .A(n305), .B(n299), .Y(n974) );
  INVX1 U791 ( .A(n974), .Y(n263) );
  AND2X1 U793 ( .A(n1508), .B(n1509), .Y(n896) );
  INVX1 U794 ( .A(n896), .Y(n264) );
  BUFX2 U797 ( .A(n897), .Y(n265) );
  INVX1 U799 ( .A(n267), .Y(n266) );
  BUFX2 U800 ( .A(n1080), .Y(n267) );
  INVX1 U803 ( .A(n1081), .Y(n268) );
  AND2X1 U804 ( .A(n720), .B(n1054), .Y(n1081) );
  INVX1 U805 ( .A(n270), .Y(n269) );
  BUFX2 U809 ( .A(n947), .Y(n270) );
  BUFX2 U810 ( .A(n1052), .Y(n271) );
  BUFX2 U812 ( .A(n1032), .Y(n272) );
  INVX1 U813 ( .A(n45), .Y(n1032) );
  INVX1 U815 ( .A(n36), .Y(n274) );
  BUFX2 U816 ( .A(n1018), .Y(n278) );
  INVX1 U818 ( .A(n46), .Y(n1018) );
  INVX1 U819 ( .A(n19), .Y(n280) );
  INVX1 U821 ( .A(n37), .Y(n281) );
  INVX1 U822 ( .A(n973), .Y(n283) );
  BUFX2 U824 ( .A(n1002), .Y(n285) );
  INVX1 U825 ( .A(n287), .Y(n286) );
  BUFX2 U827 ( .A(n866), .Y(n287) );
  OR2X1 U828 ( .A(reset), .B(n291), .Y(n816) );
  INVX1 U830 ( .A(n816), .Y(n288) );
  INVX1 U831 ( .A(n822), .Y(n289) );
  AND2X1 U833 ( .A(n962), .B(counter[0]), .Y(n1012) );
  INVX1 U834 ( .A(n1012), .Y(n290) );
  BUFX2 U836 ( .A(n837), .Y(n291) );
  INVX1 U837 ( .A(n893), .Y(n293) );
  INVX1 U839 ( .A(n42), .Y(n294) );
  INVX1 U840 ( .A(n41), .Y(n295) );
  INVX1 U842 ( .A(n895), .Y(n298) );
  BUFX2 U843 ( .A(n976), .Y(n299) );
  INVX1 U845 ( .A(n301), .Y(n300) );
  BUFX2 U846 ( .A(n1020), .Y(n301) );
  OR2X1 U848 ( .A(n461), .B(n494), .Y(n845) );
  INVX1 U849 ( .A(n845), .Y(n302) );
  INVX1 U851 ( .A(n831), .Y(n303) );
  OR2X1 U852 ( .A(n434), .B(n494), .Y(n826) );
  INVX1 U854 ( .A(n826), .Y(n304) );
  BUFX2 U855 ( .A(n975), .Y(n305) );
  INVX1 U857 ( .A(n1166), .Y(n306) );
  INVX1 U861 ( .A(n930), .Y(n307) );
  OR2X1 U862 ( .A(n365), .B(n509), .Y(n498) );
  AND2X1 U863 ( .A(n1113), .B(n1191), .Y(n1210) );
  INVX1 U864 ( .A(n1210), .Y(n308) );
  INVX1 U866 ( .A(n1439), .Y(n309) );
  BUFX2 U867 ( .A(n1150), .Y(n310) );
  BUFX2 U868 ( .A(n1151), .Y(n311) );
  INVX1 U870 ( .A(n1428), .Y(n312) );
  BUFX2 U874 ( .A(n1125), .Y(n313) );
  BUFX2 U875 ( .A(n1126), .Y(n314) );
  AND2X1 U877 ( .A(n1106), .B(n1191), .Y(n1243) );
  INVX1 U878 ( .A(n1243), .Y(n315) );
  AND2X1 U879 ( .A(state[0]), .B(n152), .Y(n732) );
  INVX1 U881 ( .A(n732), .Y(n316) );
  AND2X1 U882 ( .A(ATOMIC_cmd), .B(ATOMIC_data[15]), .Y(n1274) );
  INVX1 U883 ( .A(n1274), .Y(n317) );
  INVX1 U884 ( .A(n1438), .Y(n318) );
  BUFX2 U886 ( .A(n1148), .Y(n319) );
  BUFX2 U887 ( .A(n1149), .Y(n320) );
  INVX1 U888 ( .A(n1427), .Y(n321) );
  BUFX2 U889 ( .A(n1124), .Y(n322) );
  BUFX2 U892 ( .A(n1123), .Y(n323) );
  AND2X1 U893 ( .A(n1117), .B(n1191), .Y(n1190) );
  INVX1 U894 ( .A(n1190), .Y(n324) );
  AND2X1 U895 ( .A(n163), .B(state[0]), .Y(n776) );
  INVX1 U896 ( .A(n776), .Y(n325) );
  AND2X1 U898 ( .A(ATOMIC_cmd), .B(ATOMIC_data[14]), .Y(n1275) );
  INVX1 U899 ( .A(n1275), .Y(n326) );
  INVX1 U900 ( .A(n1436), .Y(n327) );
  BUFX2 U901 ( .A(n1141), .Y(n328) );
  BUFX2 U902 ( .A(n1142), .Y(n329) );
  INVX1 U903 ( .A(n1426), .Y(n330) );
  BUFX2 U904 ( .A(n1122), .Y(n331) );
  BUFX2 U905 ( .A(n1121), .Y(n332) );
  AND2X1 U906 ( .A(n1116), .B(n1191), .Y(n1204) );
  INVX1 U907 ( .A(n1204), .Y(n333) );
  AND2X1 U908 ( .A(n162), .B(state[0]), .Y(n772) );
  INVX1 U909 ( .A(n772), .Y(n334) );
  OR2X1 U910 ( .A(n499), .B(n462), .Y(n509) );
  AND2X1 U911 ( .A(ATOMIC_cmd), .B(ATOMIC_data[9]), .Y(n1280) );
  INVX1 U912 ( .A(n1280), .Y(n335) );
  INVX1 U913 ( .A(n1435), .Y(n336) );
  BUFX2 U914 ( .A(n1139), .Y(n337) );
  BUFX2 U915 ( .A(n1140), .Y(n338) );
  INVX1 U916 ( .A(n1425), .Y(n339) );
  BUFX2 U917 ( .A(n1119), .Y(n340) );
  BUFX2 U918 ( .A(n1118), .Y(n341) );
  AND2X1 U919 ( .A(n1111), .B(n1191), .Y(n1212) );
  INVX1 U920 ( .A(n1212), .Y(n342) );
  AND2X1 U921 ( .A(n157), .B(state[0]), .Y(n752) );
  INVX1 U922 ( .A(n752), .Y(n343) );
  AND2X1 U923 ( .A(ATOMIC_cmd), .B(ATOMIC_data[8]), .Y(n1281) );
  INVX1 U924 ( .A(n1281), .Y(n344) );
  INVX1 U925 ( .A(n1434), .Y(n345) );
  BUFX2 U926 ( .A(n1137), .Y(n346) );
  BUFX2 U927 ( .A(n1138), .Y(n347) );
  INVX1 U928 ( .A(n1424), .Y(n348) );
  BUFX2 U929 ( .A(n1105), .Y(n349) );
  BUFX2 U930 ( .A(n1104), .Y(n351) );
  AND2X1 U931 ( .A(n1110), .B(n1191), .Y(n1213) );
  INVX1 U932 ( .A(n1213), .Y(n352) );
  AND2X1 U933 ( .A(n156), .B(state[0]), .Y(n748) );
  INVX1 U934 ( .A(n748), .Y(n353) );
  AND2X1 U935 ( .A(n890), .B(n1054), .Y(n848) );
  INVX1 U936 ( .A(n848), .Y(n354) );
  AND2X1 U937 ( .A(ATOMIC_cmd), .B(ATOMIC_data[13]), .Y(n1276) );
  INVX1 U938 ( .A(n1276), .Y(n355) );
  AND2X1 U939 ( .A(ATOMIC_cmd), .B(ATOMIC_data[7]), .Y(n1282) );
  INVX1 U940 ( .A(n1282), .Y(n356) );
  INVX1 U941 ( .A(n1433), .Y(n357) );
  BUFX2 U942 ( .A(n1135), .Y(n358) );
  BUFX2 U943 ( .A(n1136), .Y(n359) );
  INVX1 U944 ( .A(n1423), .Y(n360) );
  BUFX2 U945 ( .A(n1103), .Y(n361) );
  BUFX2 U946 ( .A(n1102), .Y(n362) );
  AND2X1 U947 ( .A(n1109), .B(n1191), .Y(n1214) );
  INVX1 U948 ( .A(n1214), .Y(n363) );
  AND2X1 U949 ( .A(n155), .B(state[0]), .Y(n744) );
  INVX1 U950 ( .A(n744), .Y(n364) );
  BUFX2 U951 ( .A(n1249), .Y(n365) );
  AND2X1 U952 ( .A(n1470), .B(n432), .Y(n1184) );
  AND2X1 U953 ( .A(CMD_data_out[0]), .B(n1159), .Y(n1220) );
  INVX1 U954 ( .A(n1220), .Y(n366) );
  AND2X1 U955 ( .A(ATOMIC_cmd), .B(ATOMIC_data[12]), .Y(n1277) );
  INVX1 U956 ( .A(n1277), .Y(n367) );
  AND2X1 U957 ( .A(ATOMIC_cmd), .B(ATOMIC_data[6]), .Y(n1283) );
  INVX1 U958 ( .A(n1283), .Y(n368) );
  INVX1 U959 ( .A(n1432), .Y(n369) );
  BUFX2 U960 ( .A(n1133), .Y(n370) );
  BUFX2 U961 ( .A(n1134), .Y(n371) );
  INVX1 U962 ( .A(n1422), .Y(n372) );
  BUFX2 U963 ( .A(n1101), .Y(n373) );
  BUFX2 U964 ( .A(n1100), .Y(n374) );
  AND2X1 U965 ( .A(n1107), .B(n1191), .Y(n1217) );
  INVX1 U966 ( .A(n1217), .Y(n375) );
  AND2X1 U967 ( .A(n153), .B(state[0]), .Y(n736) );
  INVX1 U968 ( .A(n736), .Y(n376) );
  BUFX2 U969 ( .A(n1064), .Y(n377) );
  BUFX2 U970 ( .A(n1254), .Y(n378) );
  BUFX2 U971 ( .A(n844), .Y(n379) );
  OR2X1 U972 ( .A(n378), .B(n509), .Y(n728) );
  AND2X1 U973 ( .A(CMD_data_out[1]), .B(n1159), .Y(n1219) );
  INVX1 U974 ( .A(n1219), .Y(n381) );
  AND2X1 U975 ( .A(A[11]), .B(n816), .Y(n921) );
  INVX1 U976 ( .A(n921), .Y(n382) );
  AND2X1 U977 ( .A(ATOMIC_cmd), .B(ATOMIC_data[11]), .Y(n1278) );
  INVX1 U978 ( .A(n1278), .Y(n383) );
  AND2X1 U979 ( .A(ATOMIC_cmd), .B(ATOMIC_data[5]), .Y(n1284) );
  INVX1 U980 ( .A(n1284), .Y(n384) );
  INVX1 U981 ( .A(n1431), .Y(n385) );
  BUFX2 U982 ( .A(n1131), .Y(n386) );
  BUFX2 U983 ( .A(n1132), .Y(n387) );
  INVX1 U984 ( .A(n1421), .Y(n388) );
  BUFX2 U985 ( .A(n1099), .Y(n389) );
  BUFX2 U986 ( .A(n1098), .Y(n390) );
  AND2X1 U987 ( .A(n1112), .B(n1191), .Y(n1211) );
  INVX1 U988 ( .A(n1211), .Y(n391) );
  AND2X1 U989 ( .A(n158), .B(state[0]), .Y(n756) );
  INVX1 U990 ( .A(n756), .Y(n392) );
  AND2X1 U991 ( .A(n410), .B(n1054), .Y(n823) );
  INVX1 U992 ( .A(n823), .Y(n393) );
  BUFX2 U993 ( .A(n1273), .Y(n394) );
  BUFX2 U994 ( .A(n1292), .Y(n395) );
  BUFX2 U995 ( .A(n830), .Y(n396) );
  AND2X1 U996 ( .A(A[12]), .B(n816), .Y(n920) );
  INVX1 U997 ( .A(n920), .Y(n397) );
  AND2X1 U998 ( .A(ATOMIC_cmd), .B(ATOMIC_data[10]), .Y(n1279) );
  INVX1 U999 ( .A(n1279), .Y(n398) );
  AND2X1 U1000 ( .A(ATOMIC_cmd), .B(ATOMIC_data[4]), .Y(n1285) );
  INVX1 U1001 ( .A(n1285), .Y(n399) );
  INVX1 U1002 ( .A(n1430), .Y(n400) );
  BUFX2 U1003 ( .A(n1129), .Y(n401) );
  BUFX2 U1004 ( .A(n1130), .Y(n402) );
  INVX1 U1005 ( .A(n1420), .Y(n403) );
  BUFX2 U1006 ( .A(n1097), .Y(n404) );
  BUFX2 U1007 ( .A(n1096), .Y(n405) );
  AND2X1 U1008 ( .A(n1114), .B(n1191), .Y(n1208) );
  INVX1 U1009 ( .A(n1208), .Y(n406) );
  AND2X1 U1010 ( .A(n160), .B(state[0]), .Y(n764) );
  INVX1 U1011 ( .A(n764), .Y(n407) );
  AND2X1 U1012 ( .A(n962), .B(counter[4]), .Y(n1241) );
  INVX1 U1013 ( .A(n1241), .Y(n408) );
  OR2X1 U1014 ( .A(n1370), .B(n834), .Y(n1203) );
  INVX1 U1015 ( .A(n1203), .Y(n409) );
  BUFX2 U1016 ( .A(n881), .Y(n410) );
  BUFX2 U1017 ( .A(n888), .Y(n411) );
  BUFX2 U1018 ( .A(n1005), .Y(n412) );
  AND2X1 U1019 ( .A(n1061), .B(n1476), .Y(n995) );
  INVX1 U1020 ( .A(n995), .Y(n413) );
  BUFX2 U1021 ( .A(n832), .Y(n414) );
  OR2X1 U1022 ( .A(n1073), .B(n1159), .Y(n1062) );
  INVX1 U1023 ( .A(n1062), .Y(n415) );
  BUFX2 U1024 ( .A(n1076), .Y(n416) );
  AND2X1 U1025 ( .A(CMD_data_out[2]), .B(n1159), .Y(n1218) );
  INVX1 U1026 ( .A(n1218), .Y(n417) );
  AND2X1 U1027 ( .A(BA[1]), .B(n816), .Y(n919) );
  INVX1 U1028 ( .A(n919), .Y(n418) );
  AND2X1 U1029 ( .A(read_pointer[1]), .B(n712), .Y(n713) );
  INVX1 U1030 ( .A(n713), .Y(n419) );
  AND2X1 U1031 ( .A(ATOMIC_cmd), .B(ATOMIC_data[3]), .Y(n1286) );
  INVX1 U1032 ( .A(n1286), .Y(n420) );
  INVX1 U1033 ( .A(n1429), .Y(n421) );
  BUFX2 U1034 ( .A(n1127), .Y(n422) );
  BUFX2 U1035 ( .A(n1128), .Y(n423) );
  INVX1 U1036 ( .A(n1419), .Y(n424) );
  BUFX2 U1037 ( .A(n1095), .Y(n425) );
  BUFX2 U1038 ( .A(n1094), .Y(n426) );
  AND2X1 U1039 ( .A(n1108), .B(n1191), .Y(n1215) );
  INVX1 U1040 ( .A(n1215), .Y(n427) );
  AND2X1 U1041 ( .A(n154), .B(state[0]), .Y(n740) );
  INVX1 U1042 ( .A(n740), .Y(n428) );
  BUFX2 U1043 ( .A(n912), .Y(n429) );
  BUFX2 U1044 ( .A(n1238), .Y(n430) );
  BUFX2 U1045 ( .A(n1182), .Y(n431) );
  INVX1 U1046 ( .A(n1181), .Y(n432) );
  AND2X1 U1047 ( .A(n266), .B(n1476), .Y(n1027) );
  INVX1 U1048 ( .A(n1027), .Y(n433) );
  AND2X1 U1049 ( .A(n1488), .B(n1007), .Y(n969) );
  INVX1 U1050 ( .A(n969), .Y(n434) );
  BUFX2 U1051 ( .A(n1079), .Y(n435) );
  AND2X1 U1052 ( .A(BA[2]), .B(n816), .Y(n918) );
  INVX1 U1053 ( .A(n918), .Y(n436) );
  AND2X1 U1054 ( .A(ATOMIC_cmd), .B(ATOMIC_data[2]), .Y(n1287) );
  INVX1 U1055 ( .A(n1287), .Y(n437) );
  INVX1 U1056 ( .A(n1413), .Y(n438) );
  BUFX2 U1057 ( .A(n1056), .Y(n439) );
  AND2X1 U1058 ( .A(listen), .B(n1471), .Y(n1055) );
  INVX1 U1059 ( .A(n1055), .Y(n440) );
  INVX1 U1060 ( .A(n1418), .Y(n441) );
  BUFX2 U1061 ( .A(n1093), .Y(n442) );
  BUFX2 U1062 ( .A(n1092), .Y(n443) );
  INVX1 U1063 ( .A(n1466), .Y(n444) );
  AND2X1 U1064 ( .A(cas_bar), .B(n723), .Y(n1247) );
  INVX1 U1065 ( .A(n1247), .Y(n445) );
  INVX1 U1066 ( .A(n1440), .Y(n446) );
  BUFX2 U1067 ( .A(n1152), .Y(n447) );
  BUFX2 U1068 ( .A(n1153), .Y(n448) );
  BUFX2 U1069 ( .A(n1407), .Y(n449) );
  AND2X1 U1070 ( .A(n284), .B(n1472), .Y(n970) );
  INVX1 U1071 ( .A(n970), .Y(n450) );
  BUFX2 U1072 ( .A(n705), .Y(n451) );
  BUFX2 U1073 ( .A(n707), .Y(n452) );
  BUFX2 U1074 ( .A(n951), .Y(n453) );
  AND2X1 U1075 ( .A(counter[1]), .B(n1492), .Y(n958) );
  INVX1 U1076 ( .A(n958), .Y(n454) );
  AND2X1 U1077 ( .A(counter[3]), .B(n1494), .Y(n1164) );
  INVX1 U1078 ( .A(n1164), .Y(n455) );
  BUFX2 U1079 ( .A(n1242), .Y(n456) );
  AND2X1 U1080 ( .A(n1367), .B(n1364), .Y(n989) );
  INVX1 U1081 ( .A(n989), .Y(n457) );
  BUFX2 U1082 ( .A(n1240), .Y(n458) );
  BUFX2 U1083 ( .A(n500), .Y(n459) );
  AND2X1 U1084 ( .A(CMD_data_out[33]), .B(n1536), .Y(n1179) );
  INVX1 U1085 ( .A(n1179), .Y(n460) );
  BUFX2 U1086 ( .A(n829), .Y(n461) );
  BUFX2 U1087 ( .A(n1250), .Y(n462) );
  AND2X1 U1088 ( .A(n114), .B(n847), .Y(n1237) );
  INVX1 U1089 ( .A(n1237), .Y(n463) );
  AND2X1 U1090 ( .A(RETURN_address[23]), .B(reset), .Y(n729) );
  INVX1 U1091 ( .A(n729), .Y(n464) );
  AND2X1 U1092 ( .A(ATOMIC_cmd), .B(ATOMIC_data[1]), .Y(n1288) );
  INVX1 U1093 ( .A(n1288), .Y(n465) );
  INVX1 U1094 ( .A(n1465), .Y(n466) );
  AND2X1 U1095 ( .A(ras_bar), .B(n723), .Y(n1245) );
  INVX1 U1096 ( .A(n1245), .Y(n467) );
  INVX1 U1097 ( .A(n1437), .Y(n468) );
  BUFX2 U1098 ( .A(n1143), .Y(n469) );
  BUFX2 U1099 ( .A(n1145), .Y(n470) );
  INVX1 U1100 ( .A(n1416), .Y(n471) );
  BUFX2 U1101 ( .A(n1083), .Y(n472) );
  BUFX2 U1102 ( .A(n1082), .Y(n473) );
  AND2X1 U1103 ( .A(n159), .B(state[0]), .Y(n761) );
  INVX1 U1104 ( .A(n761), .Y(n474) );
  OR2X1 U1105 ( .A(n1120), .B(reset), .Y(n1234) );
  INVX1 U1106 ( .A(n1234), .Y(n475) );
  AND2X1 U1107 ( .A(n1161), .B(counter[4]), .Y(n1026) );
  INVX1 U1108 ( .A(n1026), .Y(n476) );
  BUFX2 U1109 ( .A(n709), .Y(n477) );
  AND2X1 U1110 ( .A(counter[1]), .B(counter[3]), .Y(n962) );
  INVX1 U1111 ( .A(n962), .Y(n478) );
  BUFX2 U1112 ( .A(n1258), .Y(n479) );
  INVX1 U1113 ( .A(n275), .Y(n480) );
  BUFX2 U1114 ( .A(n833), .Y(n481) );
  BUFX2 U1115 ( .A(n883), .Y(n482) );
  BUFX2 U1116 ( .A(n490), .Y(n483) );
  AND2X1 U1117 ( .A(n1494), .B(n1492), .Y(n1059) );
  INVX1 U1118 ( .A(n1059), .Y(n484) );
  AND2X1 U1119 ( .A(CMD_data_out[32]), .B(n1537), .Y(n1173) );
  INVX1 U1120 ( .A(n1173), .Y(n489) );
  OR2X1 U1121 ( .A(n266), .B(n720), .Y(n922) );
  INVX1 U1122 ( .A(n922), .Y(n494) );
  INVX1 U1123 ( .A(n435), .Y(n499) );
  AND2X1 U1124 ( .A(RETURN_address[25]), .B(reset), .Y(n811) );
  INVX1 U1125 ( .A(n811), .Y(n511) );
  AND2X1 U1126 ( .A(RETURN_address[24]), .B(reset), .Y(n809) );
  INVX1 U1127 ( .A(n809), .Y(n513) );
  AND2X1 U1128 ( .A(RETURN_address[0]), .B(reset), .Y(n807) );
  INVX1 U1129 ( .A(n807), .Y(n522) );
  AND2X1 U1130 ( .A(RETURN_address[1]), .B(reset), .Y(n805) );
  INVX1 U1131 ( .A(n805), .Y(n524) );
  AND2X1 U1132 ( .A(RETURN_address[2]), .B(reset), .Y(n803) );
  INVX1 U1133 ( .A(n803), .Y(n532) );
  AND2X1 U1134 ( .A(RETURN_address[3]), .B(reset), .Y(n775) );
  INVX1 U1135 ( .A(n775), .Y(n534) );
  AND2X1 U1136 ( .A(RETURN_address[4]), .B(reset), .Y(n773) );
  INVX1 U1137 ( .A(n773), .Y(n542) );
  AND2X1 U1138 ( .A(RETURN_address[5]), .B(reset), .Y(n771) );
  INVX1 U1139 ( .A(n771), .Y(n544) );
  AND2X1 U1140 ( .A(RETURN_address[6]), .B(reset), .Y(n769) );
  INVX1 U1141 ( .A(n769), .Y(n552) );
  AND2X1 U1142 ( .A(RETURN_address[7]), .B(reset), .Y(n767) );
  INVX1 U1143 ( .A(n767), .Y(n554) );
  AND2X1 U1144 ( .A(RETURN_address[8]), .B(reset), .Y(n765) );
  INVX1 U1145 ( .A(n765), .Y(n562) );
  AND2X1 U1146 ( .A(RETURN_address[9]), .B(reset), .Y(n757) );
  INVX1 U1147 ( .A(n757), .Y(n564) );
  AND2X1 U1148 ( .A(RETURN_address[10]), .B(reset), .Y(n755) );
  INVX1 U1149 ( .A(n755), .Y(n572) );
  AND2X1 U1150 ( .A(RETURN_address[11]), .B(reset), .Y(n753) );
  INVX1 U1151 ( .A(n753), .Y(n574) );
  AND2X1 U1152 ( .A(RETURN_address[12]), .B(reset), .Y(n751) );
  INVX1 U1153 ( .A(n751), .Y(n582) );
  AND2X1 U1154 ( .A(RETURN_address[13]), .B(reset), .Y(n749) );
  INVX1 U1155 ( .A(n749), .Y(n584) );
  AND2X1 U1156 ( .A(RETURN_address[14]), .B(reset), .Y(n747) );
  INVX1 U1157 ( .A(n747), .Y(n618) );
  AND2X1 U1158 ( .A(RETURN_address[15]), .B(reset), .Y(n745) );
  INVX1 U1159 ( .A(n745), .Y(n620) );
  AND2X1 U1160 ( .A(RETURN_address[16]), .B(reset), .Y(n743) );
  INVX1 U1161 ( .A(n743), .Y(n640) );
  AND2X1 U1162 ( .A(RETURN_address[17]), .B(reset), .Y(n741) );
  INVX1 U1163 ( .A(n741), .Y(n642) );
  AND2X1 U1164 ( .A(RETURN_address[18]), .B(reset), .Y(n739) );
  INVX1 U1165 ( .A(n739), .Y(n651) );
  AND2X1 U1166 ( .A(RETURN_address[19]), .B(reset), .Y(n737) );
  INVX1 U1167 ( .A(n737), .Y(n653) );
  AND2X1 U1168 ( .A(RETURN_address[20]), .B(reset), .Y(n735) );
  INVX1 U1169 ( .A(n735), .Y(n661) );
  AND2X1 U1170 ( .A(RETURN_address[21]), .B(reset), .Y(n733) );
  INVX1 U1171 ( .A(n733), .Y(n663) );
  AND2X1 U1172 ( .A(RETURN_address[22]), .B(reset), .Y(n731) );
  INVX1 U1173 ( .A(n731), .Y(n671) );
  AND2X1 U1174 ( .A(ATOMIC_cmd), .B(ATOMIC_data[0]), .Y(n1289) );
  INVX1 U1175 ( .A(n1289), .Y(n673) );
  AND2X1 U1176 ( .A(refresh_counter[12]), .B(n1554), .Y(n1230) );
  INVX1 U1177 ( .A(n1230), .Y(n681) );
  INVX1 U1178 ( .A(n1441), .Y(n683) );
  BUFX2 U1179 ( .A(n1155), .Y(n685) );
  BUFX2 U1180 ( .A(n1154), .Y(n686) );
  INVX1 U1181 ( .A(n1417), .Y(n687) );
  BUFX2 U1182 ( .A(n1091), .Y(n693) );
  BUFX2 U1183 ( .A(n1090), .Y(n698) );
  AND2X1 U1184 ( .A(n1115), .B(n1191), .Y(n1206) );
  INVX1 U1185 ( .A(n1206), .Y(n702) );
  AND2X1 U1186 ( .A(n161), .B(state[0]), .Y(n768) );
  INVX1 U1187 ( .A(n768), .Y(n706) );
  INVX1 U1188 ( .A(n276), .Y(n708) );
  BUFX2 U1189 ( .A(n1259), .Y(n710) );
  INVX1 U1190 ( .A(n860), .Y(n711) );
  BUFX2 U1191 ( .A(n889), .Y(n715) );
  AND2X1 U1192 ( .A(n1081), .B(n1467), .Y(n714) );
  INVX1 U1193 ( .A(n714), .Y(n716) );
  OR2X1 U1194 ( .A(n1475), .B(state[0]), .Y(n727) );
  INVX1 U1195 ( .A(n727), .Y(n720) );
  AND2X1 U1196 ( .A(n1068), .B(n1067), .Y(n1159) );
  INVX1 U1197 ( .A(n1159), .Y(n722) );
  OR2X1 U1198 ( .A(reset), .B(n1144), .Y(n1195) );
  INVX1 U1199 ( .A(n1195), .Y(n723) );
  BUFX2 U1200 ( .A(n999), .Y(n724) );
  BUFX2 U1201 ( .A(n884), .Y(n725) );
  BUFX2 U1202 ( .A(n927), .Y(n1008) );
  BUFX2 U1203 ( .A(n927), .Y(n1009) );
  BUFX2 U1204 ( .A(n926), .Y(n1003) );
  BUFX2 U1205 ( .A(n926), .Y(n1006) );
  AND2X1 U1206 ( .A(n1476), .B(n1081), .Y(n1048) );
  INVX1 U1207 ( .A(n1051), .Y(n1041) );
  INVX1 U1208 ( .A(n1051), .Y(n1040) );
  INVX1 U1209 ( .A(n1039), .Y(n1038) );
  INVX1 U1210 ( .A(reset), .Y(n1063) );
  INVX1 U1211 ( .A(reset), .Y(n1067) );
  INVX1 U1212 ( .A(n955), .Y(n1144) );
  AND2X1 U1213 ( .A(n1033), .B(n1067), .Y(n1191) );
  INVX1 U1214 ( .A(n462), .Y(n1476) );
  INVX1 U1215 ( .A(n40), .Y(n1239) );
  INVX1 U1216 ( .A(n957), .Y(n1120) );
  INVX1 U1217 ( .A(n725), .Y(n1365) );
  BUFX2 U1218 ( .A(n492), .Y(n1021) );
  INVX1 U1219 ( .A(n377), .Y(n1362) );
  BUFX2 U1220 ( .A(n492), .Y(n1024) );
  AND2X1 U1221 ( .A(n994), .B(n1067), .Y(n986) );
  BUFX2 U1222 ( .A(n515), .Y(n1036) );
  INVX1 U1223 ( .A(n479), .Y(n1360) );
  OR2X1 U1224 ( .A(n931), .B(n817), .Y(n865) );
  INVX1 U1225 ( .A(n1157), .Y(n1205) );
  INVX1 U1226 ( .A(n1085), .Y(n1051) );
  AND2X1 U1227 ( .A(n266), .B(n1157), .Y(n1085) );
  INVX1 U1228 ( .A(n1086), .Y(n1039) );
  AND2X1 U1229 ( .A(n1081), .B(n1157), .Y(n1086) );
  INVX1 U1230 ( .A(n483), .Y(n1037) );
  INVX1 U1231 ( .A(ready), .Y(n1058) );
  INVX1 U1232 ( .A(n305), .Y(n1200) );
  INVX1 U1233 ( .A(n724), .Y(n1370) );
  INVX1 U1234 ( .A(n931), .Y(n1478) );
  INVX1 U1235 ( .A(n396), .Y(n1361) );
  AND2X1 U1236 ( .A(n1483), .B(n1484), .Y(n1291) );
  INVX1 U1237 ( .A(n459), .Y(n1496) );
  AND2X1 U1238 ( .A(n1477), .B(n1371), .Y(n1260) );
  INVX1 U1239 ( .A(n1202), .Y(n1480) );
  BUFX2 U1240 ( .A(n1188), .Y(n1033) );
  AND2X1 U1241 ( .A(n1494), .B(n1371), .Y(n1007) );
  INVX1 U1242 ( .A(n950), .Y(n963) );
  INVX1 U1243 ( .A(n944), .Y(n959) );
  INVX1 U1244 ( .A(n899), .Y(n964) );
  INVX1 U1245 ( .A(n900), .Y(n967) );
  INVX1 U1246 ( .A(n902), .Y(n968) );
  INVX1 U1247 ( .A(n907), .Y(n977) );
  INVX1 U1248 ( .A(n908), .Y(n979) );
  INVX1 U1249 ( .A(n910), .Y(n981) );
  INVX1 U1250 ( .A(n911), .Y(n983) );
  INVX1 U1251 ( .A(n913), .Y(n985) );
  INVX1 U1252 ( .A(n916), .Y(n987) );
  INVX1 U1253 ( .A(n917), .Y(n990) );
  INVX1 U1254 ( .A(n925), .Y(n992) );
  INVX1 U1255 ( .A(n898), .Y(n993) );
  INVX1 U1256 ( .A(n861), .Y(n1469) );
  AND2X1 U1257 ( .A(n703), .B(n1497), .Y(n730) );
  INVX1 U1258 ( .A(n730), .Y(n501) );
  BUFX2 U1259 ( .A(n496), .Y(n1035) );
  INVX1 U1260 ( .A(n481), .Y(n1472) );
  INVX1 U1261 ( .A(n835), .Y(n1363) );
  AND2X1 U1262 ( .A(n1007), .B(n1493), .Y(n1014) );
  AND2X1 U1263 ( .A(n1491), .B(n1492), .Y(n1015) );
  AND2X1 U1264 ( .A(n688), .B(n1498), .Y(n492) );
  INVX1 U1265 ( .A(n33), .Y(n1488) );
  INVX1 U1266 ( .A(n482), .Y(n1366) );
  INVX1 U1267 ( .A(n378), .Y(n1207) );
  AND2X1 U1268 ( .A(n1161), .B(n1491), .Y(n961) );
  INVX1 U1269 ( .A(n43), .Y(n1374) );
  INVX1 U1270 ( .A(n365), .Y(n1216) );
  INVX1 U1271 ( .A(n271), .Y(n1467) );
  INVX1 U1272 ( .A(n477), .Y(n1372) );
  INVX1 U1273 ( .A(n710), .Y(n1486) );
  INVX1 U1274 ( .A(n35), .Y(n1209) );
  INVX1 U1275 ( .A(n864), .Y(n1226) );
  AND2X1 U1276 ( .A(n1068), .B(n1157), .Y(n1084) );
  INVX1 U1277 ( .A(n39), .Y(n1364) );
  INVX1 U1278 ( .A(n715), .Y(n1368) );
  INVX1 U1279 ( .A(n411), .Y(n1369) );
  INVX1 U1280 ( .A(n456), .Y(n1473) );
  INVX1 U1281 ( .A(n299), .Y(n1375) );
  INVX1 U1282 ( .A(n38), .Y(n1367) );
  INVX1 U1283 ( .A(RETURN_data[8]), .Y(n1156) );
  INVX1 U1284 ( .A(RETURN_data[13]), .Y(n1074) );
  INVX1 U1285 ( .A(RETURN_data[12]), .Y(n1075) );
  INVX1 U1286 ( .A(RETURN_data[11]), .Y(n1077) );
  INVX1 U1287 ( .A(RETURN_data[10]), .Y(n1078) );
  INVX1 U1288 ( .A(RETURN_data[9]), .Y(n1089) );
  INVX1 U1289 ( .A(RETURN_data[5]), .Y(n1178) );
  INVX1 U1290 ( .A(RETURN_data[4]), .Y(n1180) );
  INVX1 U1291 ( .A(RETURN_data[3]), .Y(n1183) );
  INVX1 U1292 ( .A(RETURN_data[2]), .Y(n1189) );
  INVX1 U1293 ( .A(RETURN_data[6]), .Y(n1172) );
  INVX1 U1294 ( .A(RETURN_data[14]), .Y(n1072) );
  INVX1 U1295 ( .A(RETURN_data[1]), .Y(n1194) );
  INVX1 U1296 ( .A(RETURN_data[7]), .Y(n1167) );
  INVX1 U1297 ( .A(RETURN_data[15]), .Y(n1070) );
  INVX1 U1298 ( .A(RETURN_data[0]), .Y(n1199) );
  AND2X1 U1299 ( .A(CMD_op[0]), .B(n703), .Y(n503) );
  AND2X1 U1300 ( .A(n688), .B(CMD_op[1]), .Y(n502) );
  AND2X1 U1301 ( .A(n1067), .B(n1498), .Y(n704) );
  AND2X1 U1302 ( .A(n1067), .B(n1499), .Y(n701) );
  INVX1 U1303 ( .A(counter[2]), .Y(n1493) );
  INVX1 U1304 ( .A(counter[0]), .Y(n1371) );
  INVX1 U1305 ( .A(counter[5]), .Y(n1489) );
  INVX1 U1306 ( .A(counter[3]), .Y(n1492) );
  INVX1 U1307 ( .A(n18), .Y(n1222) );
  INVX1 U1308 ( .A(n32), .Y(n1221) );
  INVX1 U1309 ( .A(n818), .Y(n1228) );
  AND2X1 U1310 ( .A(n961), .B(n958), .Y(n1293) );
  INVX1 U1311 ( .A(n1043), .Y(n1446) );
  INVX1 U1312 ( .A(counter[1]), .Y(n1494) );
  INVX1 U1313 ( .A(DQS_out[1]), .Y(n1502) );
  INVX1 U1314 ( .A(DQS_out[0]), .Y(n1501) );
  INVX1 U1315 ( .A(read_pointer[1]), .Y(n1533) );
  INVX1 U1316 ( .A(counter[7]), .Y(n1485) );
  INVX1 U1317 ( .A(counter[6]), .Y(n1487) );
  INVX1 U1318 ( .A(CMD_addr[23]), .Y(n1531) );
  INVX1 U1319 ( .A(CMD_addr[20]), .Y(n1528) );
  INVX1 U1320 ( .A(CMD_addr[19]), .Y(n1527) );
  INVX1 U1321 ( .A(CMD_addr[18]), .Y(n1526) );
  INVX1 U1322 ( .A(CMD_addr[17]), .Y(n1525) );
  INVX1 U1323 ( .A(CMD_addr[16]), .Y(n1524) );
  INVX1 U1324 ( .A(CMD_addr[15]), .Y(n1523) );
  INVX1 U1325 ( .A(CMD_addr[14]), .Y(n1522) );
  INVX1 U1326 ( .A(CMD_addr[13]), .Y(n1521) );
  INVX1 U1327 ( .A(CMD_addr[12]), .Y(n1520) );
  INVX1 U1328 ( .A(CMD_addr[11]), .Y(n1519) );
  INVX1 U1329 ( .A(CMD_addr[10]), .Y(n1518) );
  INVX1 U1330 ( .A(CMD_addr[9]), .Y(n1517) );
  INVX1 U1331 ( .A(CMD_addr[8]), .Y(n1516) );
  INVX1 U1332 ( .A(CMD_addr[7]), .Y(n1515) );
  INVX1 U1333 ( .A(CMD_addr[6]), .Y(n1514) );
  INVX1 U1334 ( .A(CMD_addr[5]), .Y(n1513) );
  INVX1 U1335 ( .A(CMD_addr[4]), .Y(n1512) );
  INVX1 U1336 ( .A(CMD_addr[3]), .Y(n1511) );
  INVX1 U1337 ( .A(n759), .Y(n1507) );
  INVX1 U1338 ( .A(read_pointer[0]), .Y(n1532) );
  INVX1 U1339 ( .A(counter[4]), .Y(n1491) );
  INVX1 U1340 ( .A(n394), .Y(n1490) );
  AND2X1 U1341 ( .A(n1491), .B(n1493), .Y(n1029) );
  INVX1 U1342 ( .A(DATA_data_out[15]), .Y(n1553) );
  INVX1 U1343 ( .A(DATA_data_out[0]), .Y(n1538) );
  INVX1 U1344 ( .A(n1057), .Y(n1471) );
  INVX1 U1345 ( .A(n453), .Y(n1481) );
  INVX1 U1346 ( .A(state[2]), .Y(n1475) );
  INVX1 U1347 ( .A(DATA_data_out[7]), .Y(n1545) );
  INVX1 U1348 ( .A(DATA_data_out[14]), .Y(n1552) );
  INVX1 U1349 ( .A(DATA_data_out[13]), .Y(n1551) );
  INVX1 U1350 ( .A(DATA_data_out[12]), .Y(n1550) );
  INVX1 U1351 ( .A(DATA_data_out[11]), .Y(n1549) );
  INVX1 U1352 ( .A(DATA_data_out[10]), .Y(n1548) );
  INVX1 U1353 ( .A(DATA_data_out[9]), .Y(n1547) );
  INVX1 U1354 ( .A(DATA_data_out[8]), .Y(n1546) );
  INVX1 U1355 ( .A(DATA_data_out[6]), .Y(n1544) );
  INVX1 U1356 ( .A(DATA_data_out[5]), .Y(n1543) );
  INVX1 U1357 ( .A(DATA_data_out[4]), .Y(n1542) );
  INVX1 U1358 ( .A(DATA_data_out[3]), .Y(n1541) );
  INVX1 U1359 ( .A(DATA_data_out[2]), .Y(n1540) );
  INVX1 U1360 ( .A(DATA_data_out[1]), .Y(n1539) );
  INVX1 U1361 ( .A(counter[10]), .Y(n1479) );
  AND2X1 U1362 ( .A(counter[2]), .B(n1489), .Y(n1161) );
  INVX1 U1363 ( .A(CMD_get), .Y(n1470) );
  INVX1 U1364 ( .A(DM_flag), .Y(n1510) );
  INVX1 U1365 ( .A(n34), .Y(n1482) );
  INVX1 U1366 ( .A(ck), .Y(n1554) );
  INVX1 U1367 ( .A(n31), .Y(n1251) );
  INVX1 U1368 ( .A(n30), .Y(n1252) );
  INVX1 U1369 ( .A(n21), .Y(n1358) );
  INVX1 U1370 ( .A(n22), .Y(n1357) );
  INVX1 U1371 ( .A(n23), .Y(n1290) );
  INVX1 U1372 ( .A(n24), .Y(n1272) );
  INVX1 U1373 ( .A(n25), .Y(n1269) );
  INVX1 U1374 ( .A(n26), .Y(n1267) );
  INVX1 U1375 ( .A(n27), .Y(n1262) );
  INVX1 U1376 ( .A(n28), .Y(n1261) );
  INVX1 U1377 ( .A(n29), .Y(n1255) );
  INVX1 U1378 ( .A(n20), .Y(n1359) );
  INVX1 U1379 ( .A(ATOMIC_cmd), .Y(n1053) );
  INVX1 U1380 ( .A(state[1]), .Y(n1054) );
  INVX1 U1381 ( .A(counter[11]), .Y(n1477) );
  INVX1 U1382 ( .A(counter[9]), .Y(n1483) );
  INVX1 U1383 ( .A(BLOCK_cmd), .Y(n1474) );
  INVX1 U1384 ( .A(counter[8]), .Y(n1484) );
  INVX1 U1385 ( .A(n44), .Y(n1495) );
  AND2X1 U1386 ( .A(n1067), .B(n1497), .Y(n696) );
  AND2X1 U1387 ( .A(n1488), .B(counter[6]), .Y(n1268) );
  INVX1 U1388 ( .A(CMD_sz[0]), .Y(n1503) );
  INVX1 U1389 ( .A(CMD_sz[1]), .Y(n1504) );
  INVX1 U1390 ( .A(CMD_op[0]), .Y(n1497) );
  INVX1 U1391 ( .A(CMD_data_out[31]), .Y(n1535) );
  INVX1 U1392 ( .A(state[0]), .Y(n998) );
  XOR2X1 U1393 ( .A(counter[2]), .B(n762), .Y(n905) );
  INVX1 U1394 ( .A(n762), .Y(n1509) );
  INVX1 U1395 ( .A(n760), .Y(n1508) );
  INVX1 U1396 ( .A(read_pointer[2]), .Y(n1534) );
  INVX1 U1397 ( .A(CMD_op[1]), .Y(n1498) );
  INVX1 U1398 ( .A(CMD_op[2]), .Y(n1499) );
  AND2X1 U1399 ( .A(CMD_data_out[33]), .B(CMD_data_out[32]), .Y(n1046) );
  INVX1 U1400 ( .A(CMD_addr[22]), .Y(n1530) );
  INVX1 U1401 ( .A(CMD_addr[21]), .Y(n1529) );
  INVX1 U1402 ( .A(CMD_addr[24]), .Y(n1506) );
  INVX1 U1403 ( .A(CMD_addr[25]), .Y(n1505) );
  INVX1 U1404 ( .A(refresh_counter[12]), .Y(n1468) );
  INVX1 U1405 ( .A(CMD_data_out[33]), .Y(n1537) );
  INVX1 U1406 ( .A(CMD_data_out[32]), .Y(n1536) );
  INVX1 U1407 ( .A(modify_setting), .Y(n1500) );
  MUX2X1 U1408 ( .B(n316), .A(n734), .S(state[2]), .Y(n1106) );
  MUX2X1 U1409 ( .B(n376), .A(n738), .S(state[2]), .Y(n1107) );
  MUX2X1 U1410 ( .B(n428), .A(n742), .S(state[2]), .Y(n1108) );
  MUX2X1 U1411 ( .B(n364), .A(n746), .S(state[2]), .Y(n1109) );
  MUX2X1 U1412 ( .B(n353), .A(n750), .S(state[2]), .Y(n1110) );
  MUX2X1 U1413 ( .B(n343), .A(n754), .S(state[2]), .Y(n1111) );
  MUX2X1 U1414 ( .B(n392), .A(n758), .S(state[2]), .Y(n1112) );
  MUX2X1 U1415 ( .B(n474), .A(n763), .S(state[2]), .Y(n1113) );
  MUX2X1 U1416 ( .B(n407), .A(n766), .S(state[2]), .Y(n1114) );
  MUX2X1 U1417 ( .B(n706), .A(n770), .S(state[2]), .Y(n1115) );
  MUX2X1 U1418 ( .B(n334), .A(n774), .S(state[2]), .Y(n1116) );
  MUX2X1 U1419 ( .B(n325), .A(n804), .S(state[2]), .Y(n1117) );
  MUX2X1 U1420 ( .B(n806), .A(n808), .S(state[2]), .Y(n1147) );
  MUX2X1 U1421 ( .B(n810), .A(n814), .S(state[2]), .Y(n1146) );
  MUX2X1 U1422 ( .B(n820), .A(n393), .S(state[0]), .Y(n815) );
  MUX2X1 U1423 ( .B(n1226), .A(n217), .S(state[1]), .Y(n828) );
  MUX2X1 U1424 ( .B(n843), .A(n354), .S(state[0]), .Y(n842) );
  MUX2X1 U1425 ( .B(n867), .A(n887), .S(state[0]), .Y(n862) );
  MUX2X1 U1426 ( .B(n628), .A(n152), .S(state[1]), .Y(n898) );
  MUX2X1 U1427 ( .B(n993), .A(n869), .S(state[0]), .Y(n734) );
  MUX2X1 U1428 ( .B(n629), .A(n153), .S(state[1]), .Y(n899) );
  MUX2X1 U1429 ( .B(n964), .A(n870), .S(state[0]), .Y(n738) );
  MUX2X1 U1430 ( .B(n630), .A(n154), .S(state[1]), .Y(n900) );
  MUX2X1 U1431 ( .B(n967), .A(n871), .S(state[0]), .Y(n742) );
  MUX2X1 U1432 ( .B(n631), .A(n155), .S(state[1]), .Y(n902) );
  MUX2X1 U1433 ( .B(n968), .A(n872), .S(state[0]), .Y(n746) );
  MUX2X1 U1434 ( .B(n632), .A(n156), .S(state[1]), .Y(n907) );
  MUX2X1 U1435 ( .B(n977), .A(n873), .S(state[0]), .Y(n750) );
  MUX2X1 U1436 ( .B(n633), .A(n157), .S(state[1]), .Y(n908) );
  MUX2X1 U1437 ( .B(n979), .A(n874), .S(state[0]), .Y(n754) );
  MUX2X1 U1438 ( .B(n634), .A(n158), .S(state[1]), .Y(n910) );
  MUX2X1 U1439 ( .B(n981), .A(n875), .S(state[0]), .Y(n758) );
  MUX2X1 U1440 ( .B(n635), .A(n159), .S(state[1]), .Y(n911) );
  MUX2X1 U1441 ( .B(n983), .A(n876), .S(state[0]), .Y(n763) );
  MUX2X1 U1442 ( .B(n636), .A(n160), .S(state[1]), .Y(n913) );
  MUX2X1 U1443 ( .B(n985), .A(n877), .S(state[0]), .Y(n766) );
  MUX2X1 U1444 ( .B(n637), .A(n161), .S(state[1]), .Y(n916) );
  MUX2X1 U1445 ( .B(n987), .A(n878), .S(state[0]), .Y(n770) );
  MUX2X1 U1446 ( .B(n638), .A(n162), .S(state[1]), .Y(n917) );
  MUX2X1 U1447 ( .B(n990), .A(n879), .S(state[0]), .Y(n774) );
  MUX2X1 U1448 ( .B(n639), .A(n163), .S(state[1]), .Y(n925) );
  MUX2X1 U1449 ( .B(n992), .A(n880), .S(state[0]), .Y(n804) );
  MUX2X1 U1450 ( .B(n835), .A(n835), .S(state[0]), .Y(n944) );
  MUX2X1 U1451 ( .B(n959), .A(n377), .S(state[1]), .Y(n808) );
  MUX2X1 U1452 ( .B(n708), .A(n286), .S(state[1]), .Y(n806) );
  MUX2X1 U1453 ( .B(n834), .A(n834), .S(state[0]), .Y(n950) );
  MUX2X1 U1454 ( .B(n963), .A(n1203), .S(state[1]), .Y(n814) );
  MUX2X1 U1455 ( .B(n480), .A(n286), .S(state[1]), .Y(n810) );
  MUX2X1 U1456 ( .B(n410), .A(n216), .S(state[1]), .Y(n820) );
  MUX2X1 U1457 ( .B(n212), .A(n815), .S(state[2]), .Y(n955) );
  MUX2X1 U1458 ( .B(n648), .A(n1087), .S(state[1]), .Y(n843) );
  MUX2X1 U1459 ( .B(n284), .A(n1373), .S(state[1]), .Y(n887) );
  MUX2X1 U1460 ( .B(n1469), .A(n1554), .S(state[1]), .Y(n867) );
  MUX2X1 U1461 ( .B(n862), .A(n842), .S(state[2]), .Y(n957) );
endmodule


module SSTL18DDR3DIFF ( PAD, PADN, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD,  PADN;
  wire   n1, n2, n3, n5;

  TBUFX2 b2 ( .A(A), .EN(TS), .Y(PADN) );
  TBUFX2 b1 ( .A(n5), .EN(TS), .Y(PAD) );
  NAND3X1 U2 ( .A(PAD), .B(n2), .C(RI), .Y(n1) );
  BUFX2 U1 ( .A(n1), .Y(n3) );
  INVX1 U3 ( .A(n3), .Y(Z) );
  INVX1 U4 ( .A(A), .Y(n5) );
  INVX1 U5 ( .A(PADN), .Y(n2) );
endmodule


module SSTL18DDR3_44 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_43 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_42 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_41 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_40 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_39 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_38 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_37 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_36 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_35 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n1) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_34 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n1) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_33 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n1) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_32 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n1) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_31 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n1) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_30 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_29 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n1) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_28 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n1) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_27 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n1) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_26 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_25 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n1) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_24 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_23 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n1) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_22 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n1) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_21 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n1) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_20 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n1) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_19 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n1) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_18 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n1) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_17 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n1) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_16 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n1) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_15 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n1) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_14 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n1) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_13 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n1) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_12 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n1) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_11 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n1) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_10 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n1) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_9 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n1) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_8 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n1) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_7 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n1) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_6 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n1) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_5 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  INVX1 U1 ( .A(A), .Y(n1) );
  AND2X1 U2 ( .A(RI), .B(PAD), .Y(Z) );
endmodule


module SSTL18DDR3_4 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_3 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_2 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_1 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3_0 ( PAD, Z, A, RI, TS );
  input A, RI, TS;
  output Z;
  inout PAD;
  wire   n1;

  TBUFX2 b1 ( .A(n1), .EN(TS), .Y(PAD) );
  AND2X1 U1 ( .A(RI), .B(PAD), .Y(Z) );
  INVX1 U2 ( .A(A), .Y(n1) );
endmodule


module SSTL18DDR3INTERFACE ( ck_pad, ckbar_pad, cke_pad, csbar_pad, rasbar_pad, 
        casbar_pad, webar_pad, ba_pad, a_pad, dm_pad, odt_pad, resetbar_pad, 
        dq_o, dqs_o, dqsbar_o, dq_pad, dqs_pad, dqsbar_pad, ri_i, ts_i, ck_i, 
        cke_i, csbar_i, rasbar_i, casbar_i, webar_i, ba_i, a_i, dq_i, dqs_i, 
        dqsbar_i, dm_i, odt_i, resetbar_i );
  output [2:0] ba_pad;
  output [12:0] a_pad;
  output [1:0] dm_pad;
  output [15:0] dq_o;
  output [1:0] dqs_o;
  output [1:0] dqsbar_o;
  inout [15:0] dq_pad;
  inout [1:0] dqs_pad;
  inout [1:0] dqsbar_pad;
  input [2:0] ba_i;
  input [12:0] a_i;
  input [15:0] dq_i;
  input [1:0] dqs_i;
  input [1:0] dqsbar_i;
  input [1:0] dm_i;
  input ri_i, ts_i, ck_i, cke_i, csbar_i, rasbar_i, casbar_i, webar_i, odt_i,
         resetbar_i;
  output ck_pad, ckbar_pad, cke_pad, csbar_pad, rasbar_pad, casbar_pad,
         webar_pad, odt_pad, resetbar_pad;


  SSTL18DDR3DIFF ck_sstl ( .PAD(ck_pad), .PADN(ckbar_pad), .Z(), .A(ck_i), 
        .RI(1'b0), .TS(1'b1) );
  SSTL18DDR3_44 cke_sstl ( .PAD(cke_pad), .Z(), .A(cke_i), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR3_43 casbar_sstl ( .PAD(casbar_pad), .Z(), .A(casbar_i), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_42 rasbar_sstl ( .PAD(rasbar_pad), .Z(), .A(rasbar_i), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_41 csbar_sstl ( .PAD(csbar_pad), .Z(), .A(csbar_i), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_40 webar_sstl ( .PAD(webar_pad), .Z(), .A(webar_i), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_39 odt_sstl ( .PAD(odt_pad), .Z(), .A(odt_i), .RI(1'b0), .TS(1'b1) );
  SSTL18DDR3_38 resetbar_sstl ( .PAD(resetbar_pad), .Z(), .A(resetbar_i), .RI(
        1'b0), .TS(1'b1) );
  SSTL18DDR3_37 BA_0__sstl_ba ( .PAD(ba_pad[0]), .Z(), .A(ba_i[0]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_36 BA_1__sstl_ba ( .PAD(ba_pad[1]), .Z(), .A(ba_i[1]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_35 BA_2__sstl_ba ( .PAD(ba_pad[2]), .Z(), .A(ba_i[2]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_34 A_0__sstl_a ( .PAD(a_pad[0]), .Z(), .A(a_i[0]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_33 A_1__sstl_a ( .PAD(a_pad[1]), .Z(), .A(a_i[1]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_32 A_2__sstl_a ( .PAD(a_pad[2]), .Z(), .A(a_i[2]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_31 A_3__sstl_a ( .PAD(a_pad[3]), .Z(), .A(a_i[3]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_30 A_4__sstl_a ( .PAD(a_pad[4]), .Z(), .A(a_i[4]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_29 A_5__sstl_a ( .PAD(a_pad[5]), .Z(), .A(a_i[5]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_28 A_6__sstl_a ( .PAD(a_pad[6]), .Z(), .A(a_i[6]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_27 A_7__sstl_a ( .PAD(a_pad[7]), .Z(), .A(a_i[7]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_26 A_8__sstl_a ( .PAD(a_pad[8]), .Z(), .A(a_i[8]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_25 A_9__sstl_a ( .PAD(a_pad[9]), .Z(), .A(a_i[9]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_24 A_10__sstl_a ( .PAD(a_pad[10]), .Z(), .A(a_i[10]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_23 A_11__sstl_a ( .PAD(a_pad[11]), .Z(), .A(a_i[11]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_22 A_12__sstl_a ( .PAD(a_pad[12]), .Z(), .A(a_i[12]), .RI(1'b0), 
        .TS(1'b1) );
  SSTL18DDR3_21 DQ_0__sstl_dq ( .PAD(dq_pad[0]), .Z(dq_o[0]), .A(dq_i[0]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_20 DQ_1__sstl_dq ( .PAD(dq_pad[1]), .Z(dq_o[1]), .A(dq_i[1]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_19 DQ_2__sstl_dq ( .PAD(dq_pad[2]), .Z(dq_o[2]), .A(dq_i[2]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_18 DQ_3__sstl_dq ( .PAD(dq_pad[3]), .Z(dq_o[3]), .A(dq_i[3]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_17 DQ_4__sstl_dq ( .PAD(dq_pad[4]), .Z(dq_o[4]), .A(dq_i[4]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_16 DQ_5__sstl_dq ( .PAD(dq_pad[5]), .Z(dq_o[5]), .A(dq_i[5]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_15 DQ_6__sstl_dq ( .PAD(dq_pad[6]), .Z(dq_o[6]), .A(dq_i[6]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_14 DQ_7__sstl_dq ( .PAD(dq_pad[7]), .Z(dq_o[7]), .A(dq_i[7]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_13 DQ_8__sstl_dq ( .PAD(dq_pad[8]), .Z(dq_o[8]), .A(dq_i[8]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_12 DQ_9__sstl_dq ( .PAD(dq_pad[9]), .Z(dq_o[9]), .A(dq_i[9]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_11 DQ_10__sstl_dq ( .PAD(dq_pad[10]), .Z(dq_o[10]), .A(dq_i[10]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_10 DQ_11__sstl_dq ( .PAD(dq_pad[11]), .Z(dq_o[11]), .A(dq_i[11]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_9 DQ_12__sstl_dq ( .PAD(dq_pad[12]), .Z(dq_o[12]), .A(dq_i[12]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_8 DQ_13__sstl_dq ( .PAD(dq_pad[13]), .Z(dq_o[13]), .A(dq_i[13]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_7 DQ_14__sstl_dq ( .PAD(dq_pad[14]), .Z(dq_o[14]), .A(dq_i[14]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_6 DQ_15__sstl_dq ( .PAD(dq_pad[15]), .Z(dq_o[15]), .A(dq_i[15]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_5 DQS_0__sstl_dqs ( .PAD(dqs_pad[0]), .Z(dqs_o[0]), .A(dqs_i[0]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_4 DQS_1__sstl_dqs ( .PAD(dqs_pad[1]), .Z(dqs_o[1]), .A(dqs_i[1]), 
        .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_3 DQSBAR_0__sstl_dqsbar ( .PAD(dqsbar_pad[0]), .Z(dqsbar_o[0]), 
        .A(dqsbar_i[0]), .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_2 DQSBAR_1__sstl_dqsbar ( .PAD(dqsbar_pad[1]), .Z(dqsbar_o[1]), 
        .A(dqsbar_i[1]), .RI(ri_i), .TS(ts_i) );
  SSTL18DDR3_1 DM_0__sstl_dm ( .PAD(dm_pad[0]), .Z(), .A(dm_i[0]), .RI(1'b0), 
        .TS(ts_i) );
  SSTL18DDR3_0 DM_1__sstl_dm ( .PAD(dm_pad[1]), .Z(), .A(dm_i[1]), .RI(1'b0), 
        .TS(ts_i) );
endmodule


module ddr3_controller ( dout, raddr, fillcount, validout, notfull, ready, 
        ck_pad, ckbar_pad, cke_pad, csbar_pad, rasbar_pad, casbar_pad, 
        webar_pad, ba_pad, a_pad, dm_pad, odt_pad, resetbar_pad, dq_pad, 
        dqs_pad, dqsbar_pad, clk, reset, read, cmd, sz, op, din, addr, initddr
 );
  output [15:0] dout;
  output [25:0] raddr;
  output [5:0] fillcount;
  output [2:0] ba_pad;
  output [12:0] a_pad;
  output [1:0] dm_pad;
  inout [15:0] dq_pad;
  inout [1:0] dqs_pad;
  inout [1:0] dqsbar_pad;
  input [2:0] cmd;
  input [1:0] sz;
  input [2:0] op;
  input [15:0] din;
  input [25:0] addr;
  input clk, reset, read, initddr;
  output validout, notfull, ready, ck_pad, ckbar_pad, cke_pad, csbar_pad,
         rasbar_pad, casbar_pad, webar_pad, odt_pad, resetbar_pad;
  wire   ck_i, n32, IN_put, IN_get, IN_full, CMD_get, CMD_empty, CMD_full,
         RETURN_put, RETURN_empty, RETURN_full, ready_i, init_rasbar,
         init_casbar, init_webar, init_cke, init_resetbar, rasbar, casbar,
         webar, ts_con, modify_setting, IN_BLW_put, n72, n74, n75, n76, n77,
         n78, n95, resetbar_i, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n139, n141, n142, n144, n148, n154, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n67, sub_261_A_3_, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24,
         SYNOPSYS_UNCONNECTED_25;
  wire   [15:0] IN_data_out;
  wire   [33:0] CMD_data_out;
  wire   [41:0] RETURN_data_in;
  wire   [1:0] init_ba;
  wire   [10:4] init_a;
  wire   [2:0] ba;
  wire   [12:0] a;
  wire   [1:0] dm_i;
  wire   [1:0] dqs_i;
  wire   [15:0] dq_i;
  wire   [1:0] dqs_o;
  wire   [15:0] dq_o;
  wire   [4:0] IN_BLW_counter;

  DFFPOSX1 ck_i_reg ( .D(n193), .CLK(clk), .Q(ck_i) );
  DFFPOSX1 IN_BLW_put_reg ( .D(n167), .CLK(clk), .Q(IN_BLW_put) );
  DFFPOSX1 IN_BLW_counter_reg_4_ ( .D(n166), .CLK(clk), .Q(IN_BLW_counter[4])
         );
  DFFPOSX1 IN_BLW_counter_reg_3_ ( .D(n162), .CLK(clk), .Q(IN_BLW_counter[3])
         );
  DFFPOSX1 IN_BLW_counter_reg_0_ ( .D(n165), .CLK(clk), .Q(IN_BLW_counter[0])
         );
  DFFPOSX1 IN_BLW_counter_reg_1_ ( .D(n164), .CLK(clk), .Q(IN_BLW_counter[1])
         );
  DFFPOSX1 IN_BLW_counter_reg_2_ ( .D(n163), .CLK(clk), .Q(IN_BLW_counter[2])
         );
  DFFPOSX1 validout_reg ( .D(n95), .CLK(clk), .Q(validout) );
  AOI22X1 U48 ( .A(init_webar), .B(n207), .C(webar), .D(ready_i), .Y(n119) );
  AOI22X1 U50 ( .A(init_rasbar), .B(n207), .C(rasbar), .D(ready_i), .Y(n121)
         );
  OAI21X1 U51 ( .A(n195), .B(n235), .C(n178), .Y(n162) );
  AOI22X1 U52 ( .A(n77), .B(n227), .C(sz[0]), .D(n124), .Y(n123) );
  OAI21X1 U53 ( .A(n195), .B(n212), .C(n182), .Y(n163) );
  OAI21X1 U55 ( .A(n195), .B(n236), .C(n180), .Y(n164) );
  OAI21X1 U57 ( .A(n195), .B(n74), .C(n179), .Y(n165) );
  OAI21X1 U59 ( .A(n195), .B(n234), .C(n177), .Y(n166) );
  AOI22X1 U60 ( .A(n78), .B(n227), .C(n72), .D(n124), .Y(n128) );
  NAND3X1 U62 ( .A(IN_BLW_put), .B(n191), .C(n186), .Y(n130) );
  OAI21X1 U64 ( .A(n224), .B(n188), .C(n181), .Y(n167) );
  OAI21X1 U67 ( .A(n233), .B(n191), .C(n131), .Y(n135) );
  NAND3X1 U68 ( .A(n232), .B(n231), .C(n225), .Y(n136) );
  NAND3X1 U69 ( .A(n74), .B(n236), .C(n137), .Y(n132) );
  NOR3X1 U70 ( .A(IN_BLW_counter[2]), .B(IN_BLW_counter[4]), .C(
        IN_BLW_counter[3]), .Y(n137) );
  NOR3X1 U71 ( .A(n228), .B(reset), .C(RETURN_empty), .Y(n95) );
  AOI22X1 U74 ( .A(casbar), .B(ready_i), .C(init_casbar), .D(n207), .Y(n139)
         );
  AOI22X1 U76 ( .A(ba[1]), .B(ready_i), .C(init_ba[1]), .D(n207), .Y(n141) );
  AOI22X1 U77 ( .A(ba[0]), .B(ready_i), .C(init_ba[0]), .D(n207), .Y(n142) );
  AOI22X1 U79 ( .A(a[8]), .B(ready_i), .C(init_a[8]), .D(n207), .Y(n144) );
  AOI22X1 U83 ( .A(a[4]), .B(ready_i), .C(init_a[4]), .D(n207), .Y(n148) );
  AOI22X1 U89 ( .A(a[10]), .B(ready_i), .C(init_a[10]), .D(n207), .Y(n154) );
  AOI21X1 U91 ( .A(n233), .B(n190), .C(IN_full), .Y(IN_put) );
  NAND3X1 U93 ( .A(notfull), .B(n233), .C(n159), .Y(n158) );
  OAI21X1 U94 ( .A(IN_full), .B(n229), .C(n184), .Y(n159) );
  OAI21X1 U96 ( .A(cmd[1]), .B(n230), .C(n194), .Y(n157) );
  FIFO_DEPTH_P25_WIDTH16 FIFO_IN ( .clk(clk), .reset(reset), .data_in(din), 
        .put(n189), .get(IN_get), .data_out(IN_data_out), .empty(), .full(
        IN_full), .fillcount(fillcount) );
  FIFO_DEPTH_P25_WIDTH34 FIFO_CMD ( .clk(clk), .reset(reset), .data_in({cmd, 
        addr, sz, op}), .put(n225), .get(CMD_get), .data_out(CMD_data_out), 
        .empty(CMD_empty), .full(CMD_full), .fillcount({SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6}) );
  FIFO_DEPTH_P25_WIDTH42 FIFO_RETURN ( .clk(clk), .reset(reset), .data_in(
        RETURN_data_in), .put(RETURN_put), .get(read), .data_out({raddr, dout}), .empty(RETURN_empty), .full(RETURN_full), .fillcount({SYNOPSYS_UNCONNECTED_7, 
        SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12}) );
  ddr3_init_engine XINIT ( .ready(ready_i), .csbar(), .rasbar(init_rasbar), 
        .casbar(init_casbar), .webar(init_webar), .ba({SYNOPSYS_UNCONNECTED_13, 
        init_ba}), .a({SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        init_a[10], SYNOPSYS_UNCONNECTED_16, init_a[8], 
        SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, 
        SYNOPSYS_UNCONNECTED_19, init_a[4], SYNOPSYS_UNCONNECTED_20, 
        SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22, 
        SYNOPSYS_UNCONNECTED_23}), .odt(), .ts_con(), .cke(init_cke), 
        .resetbar(init_resetbar), .clk(clk), .reset(reset), .init(initddr), 
        .ck(ck_i) );
  Processing_logic XPL ( .DATA_get(IN_get), .CMD_get(CMD_get), .RETURN_put(
        RETURN_put), .RETURN_address(RETURN_data_in[41:16]), .RETURN_data(
        RETURN_data_in[15:0]), .cs_bar(), .ras_bar(rasbar), .cas_bar(casbar), 
        .we_bar(webar), .BA(ba), .A(a), .DM(dm_i), .DQS_out(dqs_i), .DQ_out(
        dq_i), .ts_con(ts_con), .modify_setting(modify_setting), .clk(clk), 
        .ck(ck_i), .reset(reset), .ready(ready_i), .CMD_empty(CMD_empty), 
        .CMD_data_out(CMD_data_out), .DATA_data_out(IN_data_out), 
        .RETURN_full(RETURN_full), .DQS_in(dqs_o), .DQ_in(dq_o) );
  SSTL18DDR3INTERFACE XSSTL ( .ck_pad(ck_pad), .ckbar_pad(ckbar_pad), 
        .cke_pad(cke_pad), .csbar_pad(csbar_pad), .rasbar_pad(rasbar_pad), 
        .casbar_pad(casbar_pad), .webar_pad(webar_pad), .ba_pad(ba_pad), 
        .a_pad(a_pad), .dm_pad(dm_pad), .odt_pad(odt_pad), .resetbar_pad(
        resetbar_pad), .dq_o(dq_o), .dqs_o(dqs_o), .dqsbar_o({
        SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25}), .dq_pad(dq_pad), 
        .dqs_pad(dqs_pad), .dqsbar_pad(dqsbar_pad), .ri_i(1'b1), .ts_i(n120), 
        .ck_i(ck_i), .cke_i(init_cke), .csbar_i(1'b0), .rasbar_i(n215), 
        .casbar_i(n214), .webar_i(n218), .ba_i({n196, n223, n222}), .a_i({n206, 
        n205, n221, n204, n220, n203, n202, n201, n219, n200, n199, n198, n197}), .dq_i(dq_i), .dqs_i(dqs_i), .dqsbar_i({n217, n216}), .dm_i(dm_i), .odt_i(
        1'b0), .resetbar_i(resetbar_i) );
  AND2X1 U98 ( .A(n208), .B(n176), .Y(n131) );
  AND2X1 U99 ( .A(n131), .B(n185), .Y(n122) );
  OR2X1 U100 ( .A(n192), .B(IN_BLW_counter[3]), .Y(n211) );
  BUFX2 U101 ( .A(n154), .Y(n168) );
  BUFX2 U102 ( .A(n148), .Y(n169) );
  BUFX2 U103 ( .A(n144), .Y(n170) );
  BUFX2 U104 ( .A(n142), .Y(n171) );
  BUFX2 U105 ( .A(n141), .Y(n172) );
  BUFX2 U106 ( .A(n139), .Y(n173) );
  BUFX2 U107 ( .A(n121), .Y(n174) );
  BUFX2 U108 ( .A(n119), .Y(n175) );
  BUFX2 U109 ( .A(n136), .Y(n176) );
  BUFX2 U110 ( .A(n128), .Y(n177) );
  BUFX2 U111 ( .A(n123), .Y(n178) );
  AND2X1 U112 ( .A(n74), .B(n227), .Y(n127) );
  INVX1 U113 ( .A(n127), .Y(n179) );
  BUFX2 U114 ( .A(n126), .Y(n180) );
  AND2X1 U115 ( .A(n224), .B(IN_BLW_put), .Y(n134) );
  INVX1 U116 ( .A(n134), .Y(n181) );
  BUFX2 U117 ( .A(n125), .Y(n182) );
  AND2X1 U118 ( .A(n129), .B(n195), .Y(n124) );
  BUFX2 U119 ( .A(n158), .Y(n183) );
  AND2X1 U120 ( .A(cmd[0]), .B(n230), .Y(n160) );
  INVX1 U121 ( .A(n160), .Y(n184) );
  BUFX2 U122 ( .A(n130), .Y(n185) );
  OR2X1 U123 ( .A(reset), .B(IN_full), .Y(n133) );
  INVX1 U124 ( .A(n133), .Y(n186) );
  AND2X1 U125 ( .A(n236), .B(n74), .Y(n209) );
  INVX1 U126 ( .A(n209), .Y(n187) );
  AND2X1 U127 ( .A(n233), .B(n208), .Y(n129) );
  INVX1 U128 ( .A(n129), .Y(n188) );
  BUFX2 U129 ( .A(IN_put), .Y(n189) );
  AND2X1 U130 ( .A(n157), .B(notfull), .Y(n156) );
  INVX1 U131 ( .A(n156), .Y(n190) );
  BUFX2 U132 ( .A(n132), .Y(n191) );
  AND2X1 U133 ( .A(n209), .B(n212), .Y(n210) );
  INVX1 U134 ( .A(n210), .Y(n192) );
  AND2X1 U135 ( .A(ts_con), .B(ready_i), .Y(n120) );
  OR2X1 U136 ( .A(reset), .B(ck_i), .Y(n32) );
  INVX1 U137 ( .A(n32), .Y(n193) );
  AND2X1 U138 ( .A(cmd[1]), .B(n232), .Y(n161) );
  INVX1 U139 ( .A(n161), .Y(n194) );
  INVX1 U140 ( .A(n122), .Y(n195) );
  INVX1 U141 ( .A(n185), .Y(n227) );
  INVX1 U142 ( .A(n157), .Y(n229) );
  INVX1 U143 ( .A(read), .Y(n228) );
  INVX1 U144 ( .A(n135), .Y(n224) );
  INVX1 U145 ( .A(n183), .Y(n225) );
  INVX1 U146 ( .A(IN_BLW_counter[3]), .Y(n235) );
  INVX1 U147 ( .A(IN_BLW_counter[4]), .Y(n234) );
  INVX1 U148 ( .A(cmd[1]), .Y(n231) );
  INVX1 U149 ( .A(ready_i), .Y(n207) );
  INVX1 U150 ( .A(IN_BLW_put), .Y(n233) );
  INVX1 U151 ( .A(CMD_full), .Y(notfull) );
  AND2X1 U152 ( .A(init_resetbar), .B(n208), .Y(resetbar_i) );
  INVX1 U153 ( .A(sz[0]), .Y(sub_261_A_3_) );
  INVX1 U154 ( .A(reset), .Y(n208) );
  INVX1 U155 ( .A(cmd[2]), .Y(n230) );
  INVX1 U156 ( .A(cmd[0]), .Y(n232) );
  INVX1 U157 ( .A(IN_BLW_counter[0]), .Y(n74) );
  INVX1 U158 ( .A(IN_BLW_counter[2]), .Y(n212) );
  INVX1 U159 ( .A(IN_BLW_counter[1]), .Y(n236) );
  INVX1 U160 ( .A(n174), .Y(n215) );
  INVX1 U161 ( .A(n175), .Y(n218) );
  INVX1 U162 ( .A(n173), .Y(n214) );
  INVX1 U163 ( .A(n171), .Y(n222) );
  INVX1 U164 ( .A(n172), .Y(n223) );
  INVX1 U165 ( .A(n169), .Y(n219) );
  INVX1 U166 ( .A(n170), .Y(n220) );
  INVX1 U167 ( .A(n168), .Y(n221) );
  AND2X1 U168 ( .A(modify_setting), .B(ready_i), .Y(ready) );
  INVX1 U169 ( .A(dqs_i[0]), .Y(n216) );
  INVX1 U170 ( .A(dqs_i[1]), .Y(n217) );
  AND2X1 U171 ( .A(ba[2]), .B(ready_i), .Y(n196) );
  AND2X1 U172 ( .A(a[0]), .B(ready_i), .Y(n197) );
  AND2X1 U173 ( .A(a[1]), .B(ready_i), .Y(n198) );
  AND2X1 U174 ( .A(a[2]), .B(ready_i), .Y(n199) );
  AND2X1 U175 ( .A(a[3]), .B(ready_i), .Y(n200) );
  AND2X1 U176 ( .A(a[5]), .B(ready_i), .Y(n201) );
  AND2X1 U177 ( .A(a[6]), .B(ready_i), .Y(n202) );
  AND2X1 U178 ( .A(a[7]), .B(ready_i), .Y(n203) );
  AND2X1 U179 ( .A(a[9]), .B(ready_i), .Y(n204) );
  AND2X1 U180 ( .A(a[11]), .B(ready_i), .Y(n205) );
  AND2X1 U181 ( .A(a[12]), .B(ready_i), .Y(n206) );
  XNOR2X1 U182 ( .A(n67), .B(sub_261_A_3_), .Y(n72) );
  OAI21X1 U183 ( .A(n74), .B(n236), .C(n187), .Y(n75) );
  OAI21X1 U184 ( .A(n209), .B(n212), .C(n192), .Y(n76) );
  XNOR2X1 U185 ( .A(IN_BLW_counter[3]), .B(n192), .Y(n77) );
  XNOR2X1 U186 ( .A(IN_BLW_counter[4]), .B(n211), .Y(n78) );
  AOI21X1 U189 ( .A(n76), .B(n227), .C(n124), .Y(n125) );
  AOI21X1 U190 ( .A(n75), .B(n227), .C(n124), .Y(n126) );
  XOR2X1 U191 ( .A(sz[1]), .B(sz[0]), .Y(n67) );
endmodule

