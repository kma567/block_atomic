/////////////////////////////////////////////////////////////////////
// 
// Filename        : ddr2_ring_buffer.v
// Description     : DDR2 8 deep input ring buffer 
//                   Strobe filter and a delay line for strobe
// Author          : Rashed Bhatti
// Modified	       : Tzu-Ching Lin
/////////////////////////////////////////////////////////////////////
`timescale 1ns/10ps


module ddr3_ring_buffer8 (dout, listen, strobe, readPtr, din, reset);
   input listen;   // A cycle long pulse after which ring buffer would start paying attention towards the incoming strobe
   input [1:0] strobe;   // After listen the ring buffer would capture 4 data at every edges of strobe
   input reset;
   input [15:0]  din;
   input [2:0] 	 readPtr; // Read pointer, the contol logic should provide the read pointer
   output [15:0] dout;
 
   reg 	[15:0] 	dout;   
   reg 	[15:0] 	r0, r1, r2, r3, r4, r5, r6, r7;
   reg 			F0;
   wire 		fStrobe, fStrobeBar;
   wire	[3:0]	pStrobe, nStrobe;
   wire			dStrobe0, dStrobe1, dStrobe2, dStrobe3, dStrobe4, dStrobe5, dnStrobe, dpStrobe;
   reg 	[1:0] 	count;

// Delayline for strobe   
// --------------------
// To tell the sysnopsys not to remove the following delay cells 
// use the following line in constraint file
// set_dont_touch [ find cell DELAY*]
// get_attribute [ find cell DELAY*] dont_touch
    CLKBUF2 DELAY0 (.Y(dStrobe0), .A(strobe[1] & F0));
    CLKBUF2 DELAY1 (.Y(dStrobe1), .A(dStrobe0)); 
    CLKBUF2 DELAY2 (.Y(dStrobe2), .A(dStrobe1));
	CLKBUF2 DELAY3 (.Y(dnStrobe), .A(dStrobe2));
    
	CLKBUF2 DELAYN0 (.Y(nStrobe[0]), .A(dnStrobe));
	CLKBUF2 DELAYN1 (.Y(nStrobe[1]), .A(dnStrobe));
	CLKBUF2 DELAYN2 (.Y(nStrobe[2]), .A(dnStrobe));
	CLKBUF2 DELAYN3 (.Y(nStrobe[3]), .A(dnStrobe));
	
	CLKBUF2 DELAY4 (.Y(dStrobe3),  .A(strobe[0] & F0));
	CLKBUF2 DELAY5 (.Y(dStrobe4),  .A(dStrobe3));
	CLKBUF2 DELAY6 (.Y(dStrobe5),  .A(dStrobe4));
	CLKBUF2 DELAY7 (.Y(dpStrobe),  .A(dStrobe5));
	
	CLKBUF2 DELAYP0 (.Y(pStrobe[0]), .A(dpStrobe));
	CLKBUF2 DELAYP1 (.Y(pStrobe[1]), .A(dpStrobe));
	CLKBUF2 DELAYP2 (.Y(pStrobe[2]), .A(dpStrobe));
	CLKBUF2 DELAYP3 (.Y(pStrobe[3]), .A(dpStrobe));
	
	
	
// strobe filter
// -------------   
//     strobe   XXXX___________/-----\_____/-----\_____/-----\_____/-----\______XXXXX
//	  
//     listen   _____/-----\______________________________________________________
//	  
//     F0       ______/----------------------------------------------------\________
//   
//     fStrobe  __________________/-----\_____/-----\_____/-----\_____/-----\________
//
//     count    -----0000000000000000000011111111111122222222222233333333333300000000



   always @(posedge fStrobeBar, posedge listen, posedge reset)
   begin
		if (reset)
		begin			 
			F0 <= 0;
			count <= 0;
		end
		else if (listen)
			F0 <= 1;
		else
		begin
			if (count < 3)
				count <= count + 1;
			else if (count == 3)
			begin
				count <= 0;
				F0 <= 0;
			end
		end // else: !if(listen)
	end // always @ (posedge fStrobeBar or posedge listen or posedge reset)
   
   //assign fStrobe = Strobe & F0;
   //assign pStrobe = strobe[0] & F0;
   //assign nStrobe = dStrobe1 & F0;
   assign fStrobeBar = ~dStrobe0;


// Capture data at the edges
// -------------------------  
/*    always @(posedge pStrobe)
	 case (count)
	   0: r0 <= din;   
	   1: r2 <= din;
	   2: r4 <= din;
	   3: r6 <= din;
	 endcase // case(counter)
   always @(negedge nStrobe)
	 case (count)
	   0: r1 <= din;   
	   1: r3 <= din;
	   2: r5 <= din;
	   3: r7 <= din;
	 endcase // case(counter) */
	 
	always @(posedge pStrobe[0])
	begin
		if (count == 0)
			r0 <= din;
	end
	
	always @(posedge pStrobe[1])
	begin
		if (count == 1)
			r2 <= din;
	end
	
	always @(posedge pStrobe[2])
	begin
		if (count == 2)
			r4 <= din;
	end
	
	always @(posedge pStrobe[3])
	begin
		if (count == 3)
			r6 <= din;
	end
	
	always @(negedge nStrobe[0])
	begin
		if (count == 0)
			r1 <= din;
	end
	
	always @(negedge nStrobe[1])
	begin
		if (count == 1)
			r3 <= din;
	end
	
	always @(negedge nStrobe[2])
	begin
		if (count == 2)
			r5 <= din;
	end
	
	always @(negedge nStrobe[3])
	begin
		if (count == 3)
			r7 <= din;
	end


// Read data
// ---------
   always @ (r0 or r1 or r2 or r3 or r4 or r5 or r6 or r7 or readPtr)
	 begin
		case (readPtr) 
		  3'b000: dout = r0;
		  3'b001: dout = r1;
		  3'b010: dout = r2;
		  3'b011: dout = r3;
		  3'b100: dout = r4;
		  3'b101: dout = r5;
		  3'b110: dout = r6;
		  3'b111: dout = r7;
		  default: dout = r0;
		endcase // case (readPtr)
	 end // always (r0 or r1 or r2 or r3 or r4 or readPtr)
   
   
endmodule // ddr2_ring_buffer8
